
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity PCIe_UserLogic_00 is
  port (
    bram_rd_dout        : in  std_logic_vector(63 downto 0);
    debug_in_1i         : in  std_logic_vector(31 downto 0);
    debug_in_2i         : in  std_logic_vector(31 downto 0);
    debug_in_3i         : in  std_logic_vector(31 downto 0);
    debug_in_4i         : in  std_logic_vector(31 downto 0);
    dma_host2board_busy : in  std_logic;
    dma_host2board_done : in  std_logic;
    fifo_rd_count       : in  std_logic_vector(14 downto 0);
    fifo_rd_dout        : in  std_logic_vector(71 downto 0);
    fifo_rd_empty       : in  std_logic;
    fifo_rd_pempty      : in  std_logic;
    fifo_rd_valid       : in  std_logic;
    fifo_wr_count       : in  std_logic_vector(14 downto 0);
    fifo_wr_full        : in  std_logic;
    fifo_wr_pfull       : in  std_logic;
    inout_logic_cw_ce   : in  std_logic := '1';
    inout_logic_cw_clk  : in  std_logic;
    reg01_td            : in  std_logic_vector(31 downto 0);
    reg01_tv            : in  std_logic;
    reg02_td            : in  std_logic_vector(31 downto 0);
    reg02_tv            : in  std_logic;
    reg03_td            : in  std_logic_vector(31 downto 0);
    reg03_tv            : in  std_logic;
    reg04_td            : in  std_logic_vector(31 downto 0);
    reg04_tv            : in  std_logic;
    reg05_td            : in  std_logic_vector(31 downto 0);
    reg05_tv            : in  std_logic;
    reg06_td            : in  std_logic_vector(31 downto 0);
    reg06_tv            : in  std_logic;
    reg07_td            : in  std_logic_vector(31 downto 0);
    reg07_tv            : in  std_logic;
    reg08_td            : in  std_logic_vector(31 downto 0);
    reg08_tv            : in  std_logic;
    reg09_td            : in  std_logic_vector(31 downto 0);
    reg09_tv            : in  std_logic;
    reg10_td            : in  std_logic_vector(31 downto 0);
    reg10_tv            : in  std_logic;
    reg11_td            : in  std_logic_vector(31 downto 0);
    reg11_tv            : in  std_logic;
    reg12_td            : in  std_logic_vector(31 downto 0);
    reg12_tv            : in  std_logic;
    reg13_td            : in  std_logic_vector(31 downto 0);
    reg13_tv            : in  std_logic;
    reg14_td            : in  std_logic_vector(31 downto 0);
    reg14_tv            : in  std_logic;
    rst_i               : in  std_logic;
    user_logic_cw_ce    : in  std_logic := '1';
    user_logic_cw_clk   : in  std_logic;
    bram_rd_addr        : out std_logic_vector(11 downto 0);
    bram_wr_addr        : out std_logic_vector(11 downto 0);
    bram_wr_din         : out std_logic_vector(63 downto 0);
    bram_wr_en          : out std_logic_vector(7 downto 0);
    fifo_rd_en          : out std_logic;
    fifo_wr_din         : out std_logic_vector(71 downto 0);
    fifo_wr_en          : out std_logic;
    reg01_rd            : out std_logic_vector(31 downto 0);
    reg01_rv            : out std_logic;
    reg02_rd            : out std_logic_vector(31 downto 0);
    reg02_rv            : out std_logic;
    reg03_rd            : out std_logic_vector(31 downto 0);
    reg03_rv            : out std_logic;
    reg04_rd            : out std_logic_vector(31 downto 0);
    reg04_rv            : out std_logic;
    reg05_rd            : out std_logic_vector(31 downto 0);
    reg05_rv            : out std_logic;
    reg06_rd            : out std_logic_vector(31 downto 0);
    reg06_rv            : out std_logic;
    reg07_rd            : out std_logic_vector(31 downto 0);
    reg07_rv            : out std_logic;
    reg08_rd            : out std_logic_vector(31 downto 0);
    reg08_rv            : out std_logic;
    reg09_rd            : out std_logic_vector(31 downto 0);
    reg09_rv            : out std_logic;
    reg10_rd            : out std_logic_vector(31 downto 0);
    reg10_rv            : out std_logic;
    reg11_rd            : out std_logic_vector(31 downto 0);
    reg11_rv            : out std_logic;
    reg12_rd            : out std_logic_vector(31 downto 0);
    reg12_rv            : out std_logic;
    reg13_rd            : out std_logic_vector(31 downto 0);
    reg13_rv            : out std_logic;
    reg14_rd            : out std_logic_vector(31 downto 0);
    reg14_rv            : out std_logic;
    rst_o               : out std_logic;
    user_int_1o         : out std_logic;
    user_int_2o         : out std_logic;
    user_int_3o         : out std_logic
    );
end PCIe_UserLogic_00;

architecture structural of PCIe_UserLogic_00 is

begin
  
  bram_rd_addr <= (others => '0');
  bram_wr_addr <= (others => '0');
  bram_wr_din  <= (others => '0');
  bram_wr_en   <= (others => '0');
  fifo_rd_en   <= '0';
  fifo_wr_din  <= (others => '0');
  fifo_wr_en   <= '0';
  reg01_rd     <= (others => '0');
  reg01_rv     <= '0';
  reg02_rd     <= (others => '0');
  reg02_rv     <= '0';
  reg03_rd     <= (others => '0');
  reg03_rv     <= '0';
  reg04_rd     <= (others => '0');
  reg04_rv     <= '0';
  reg05_rd     <= (others => '0');
  reg05_rv     <= '0';
  reg06_rd     <= (others => '0');
  reg06_rv     <= '0';
  reg07_rd     <= (others => '0');
  reg07_rv     <= '0';
  reg08_rd     <= (others => '0');
  reg08_rv     <= '0';
  reg09_rd     <= (others => '0');
  reg09_rv     <= '0';
  reg10_rd     <= (others => '0');
  reg10_rv     <= '0';
  reg11_rd     <= (others => '0');
  reg11_rv     <= '0';
  reg12_rd     <= (others => '0');
  reg12_rv     <= '0';
  reg13_rd     <= (others => '0');
  reg13_rv     <= '0';
  reg14_rd     <= (others => '0');
  reg14_rv     <= '0';
  rst_o        <= '0';
  user_int_1o  <= '0';
  user_int_2o  <= '0';
  user_int_3o  <= '0';

end structural;
