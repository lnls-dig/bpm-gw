`define ADDR_ORBIT_INTLK_CTRL          6'h0
`define ORBIT_INTLK_CTRL_EN_OFFSET 0
`define ORBIT_INTLK_CTRL_EN 32'h00000001
`define ORBIT_INTLK_CTRL_CLR_OFFSET 1
`define ORBIT_INTLK_CTRL_CLR 32'h00000002
`define ORBIT_INTLK_CTRL_MIN_SUM_EN_OFFSET 2
`define ORBIT_INTLK_CTRL_MIN_SUM_EN 32'h00000004
`define ORBIT_INTLK_CTRL_TRANS_EN_OFFSET 3
`define ORBIT_INTLK_CTRL_TRANS_EN 32'h00000008
`define ORBIT_INTLK_CTRL_TRANS_CLR_OFFSET 4
`define ORBIT_INTLK_CTRL_TRANS_CLR 32'h00000010
`define ORBIT_INTLK_CTRL_ANG_EN_OFFSET 5
`define ORBIT_INTLK_CTRL_ANG_EN 32'h00000020
`define ORBIT_INTLK_CTRL_ANG_CLR_OFFSET 6
`define ORBIT_INTLK_CTRL_ANG_CLR 32'h00000040
`define ORBIT_INTLK_CTRL_RESERVED_OFFSET 7
`define ORBIT_INTLK_CTRL_RESERVED 32'h7fffff80
`define ADDR_ORBIT_INTLK_STS           6'h4
`define ORBIT_INTLK_STS_TRANS_BIGGER_X_OFFSET 0
`define ORBIT_INTLK_STS_TRANS_BIGGER_X 32'h00000001
`define ORBIT_INTLK_STS_TRANS_BIGGER_Y_OFFSET 1
`define ORBIT_INTLK_STS_TRANS_BIGGER_Y 32'h00000002
`define ORBIT_INTLK_STS_TRANS_BIGGER_LTC_X_OFFSET 2
`define ORBIT_INTLK_STS_TRANS_BIGGER_LTC_X 32'h00000004
`define ORBIT_INTLK_STS_TRANS_BIGGER_LTC_Y_OFFSET 3
`define ORBIT_INTLK_STS_TRANS_BIGGER_LTC_Y 32'h00000008
`define ORBIT_INTLK_STS_TRANS_BIGGER_ANY_OFFSET 4
`define ORBIT_INTLK_STS_TRANS_BIGGER_ANY 32'h00000010
`define ORBIT_INTLK_STS_TRANS_BIGGER_OFFSET 5
`define ORBIT_INTLK_STS_TRANS_BIGGER 32'h00000020
`define ORBIT_INTLK_STS_TRANS_BIGGER_LTC_OFFSET 6
`define ORBIT_INTLK_STS_TRANS_BIGGER_LTC 32'h00000040
`define ORBIT_INTLK_STS_ANG_BIGGER_X_OFFSET 7
`define ORBIT_INTLK_STS_ANG_BIGGER_X 32'h00000080
`define ORBIT_INTLK_STS_ANG_BIGGER_Y_OFFSET 8
`define ORBIT_INTLK_STS_ANG_BIGGER_Y 32'h00000100
`define ORBIT_INTLK_STS_ANG_BIGGER_LTC_X_OFFSET 9
`define ORBIT_INTLK_STS_ANG_BIGGER_LTC_X 32'h00000200
`define ORBIT_INTLK_STS_ANG_BIGGER_LTC_Y_OFFSET 10
`define ORBIT_INTLK_STS_ANG_BIGGER_LTC_Y 32'h00000400
`define ORBIT_INTLK_STS_ANG_BIGGER_ANY_OFFSET 11
`define ORBIT_INTLK_STS_ANG_BIGGER_ANY 32'h00000800
`define ORBIT_INTLK_STS_ANG_BIGGER_OFFSET 12
`define ORBIT_INTLK_STS_ANG_BIGGER 32'h00001000
`define ORBIT_INTLK_STS_ANG_BIGGER_LTC_OFFSET 13
`define ORBIT_INTLK_STS_ANG_BIGGER_LTC 32'h00002000
`define ORBIT_INTLK_STS_INTLK_BIGGER_OFFSET 14
`define ORBIT_INTLK_STS_INTLK_BIGGER 32'h00004000
`define ORBIT_INTLK_STS_INTLK_BIGGER_LTC_OFFSET 15
`define ORBIT_INTLK_STS_INTLK_BIGGER_LTC 32'h00008000
`define ORBIT_INTLK_STS_TRANS_SMALLER_X_OFFSET 16
`define ORBIT_INTLK_STS_TRANS_SMALLER_X 32'h00010000
`define ORBIT_INTLK_STS_TRANS_SMALLER_Y_OFFSET 17
`define ORBIT_INTLK_STS_TRANS_SMALLER_Y 32'h00020000
`define ORBIT_INTLK_STS_TRANS_SMALLER_LTC_X_OFFSET 18
`define ORBIT_INTLK_STS_TRANS_SMALLER_LTC_X 32'h00040000
`define ORBIT_INTLK_STS_TRANS_SMALLER_LTC_Y_OFFSET 19
`define ORBIT_INTLK_STS_TRANS_SMALLER_LTC_Y 32'h00080000
`define ORBIT_INTLK_STS_TRANS_SMALLER_ANY_OFFSET 20
`define ORBIT_INTLK_STS_TRANS_SMALLER_ANY 32'h00100000
`define ORBIT_INTLK_STS_TRANS_SMALLER_OFFSET 21
`define ORBIT_INTLK_STS_TRANS_SMALLER 32'h00200000
`define ORBIT_INTLK_STS_TRANS_SMALLER_LTC_OFFSET 22
`define ORBIT_INTLK_STS_TRANS_SMALLER_LTC 32'h00400000
`define ORBIT_INTLK_STS_ANG_SMALLER_X_OFFSET 23
`define ORBIT_INTLK_STS_ANG_SMALLER_X 32'h00800000
`define ORBIT_INTLK_STS_ANG_SMALLER_Y_OFFSET 24
`define ORBIT_INTLK_STS_ANG_SMALLER_Y 32'h01000000
`define ORBIT_INTLK_STS_ANG_SMALLER_LTC_X_OFFSET 25
`define ORBIT_INTLK_STS_ANG_SMALLER_LTC_X 32'h02000000
`define ORBIT_INTLK_STS_ANG_SMALLER_LTC_Y_OFFSET 26
`define ORBIT_INTLK_STS_ANG_SMALLER_LTC_Y 32'h04000000
`define ORBIT_INTLK_STS_ANG_SMALLER_ANY_OFFSET 27
`define ORBIT_INTLK_STS_ANG_SMALLER_ANY 32'h08000000
`define ORBIT_INTLK_STS_ANG_SMALLER_OFFSET 28
`define ORBIT_INTLK_STS_ANG_SMALLER 32'h10000000
`define ORBIT_INTLK_STS_ANG_SMALLER_LTC_OFFSET 29
`define ORBIT_INTLK_STS_ANG_SMALLER_LTC 32'h20000000
`define ORBIT_INTLK_STS_RESERVED_OFFSET 30
`define ORBIT_INTLK_STS_RESERVED 32'hc0000000
`define ADDR_ORBIT_INTLK_MIN_SUM       6'h8
`define ADDR_ORBIT_INTLK_TRANS_MAX_X   6'hc
`define ADDR_ORBIT_INTLK_TRANS_MAX_Y   6'h10
`define ADDR_ORBIT_INTLK_ANG_MAX_X     6'h14
`define ADDR_ORBIT_INTLK_ANG_MAX_Y     6'h18
`define ADDR_ORBIT_INTLK_TRANS_MIN_X   6'h1c
`define ADDR_ORBIT_INTLK_TRANS_MIN_Y   6'h20
`define ADDR_ORBIT_INTLK_ANG_MIN_X     6'h24
`define ADDR_ORBIT_INTLK_ANG_MIN_Y     6'h28
