`define ADDR_ACQ_CORE_CTL              8'h0
`define ACQ_CORE_CTL_FSM_START_ACQ_OFFSET 0
`define ACQ_CORE_CTL_FSM_START_ACQ 32'h00000001
`define ACQ_CORE_CTL_FSM_STOP_ACQ_OFFSET 1
`define ACQ_CORE_CTL_FSM_STOP_ACQ 32'h00000002
`define ACQ_CORE_CTL_RESERVED1_OFFSET 2
`define ACQ_CORE_CTL_RESERVED1 32'h0000fffc
`define ACQ_CORE_CTL_FSM_ACQ_NOW_OFFSET 16
`define ACQ_CORE_CTL_FSM_ACQ_NOW 32'h00010000
`define ACQ_CORE_CTL_RESERVED2_OFFSET 17
`define ACQ_CORE_CTL_RESERVED2 32'hfffe0000
`define ADDR_ACQ_CORE_STA              8'h4
`define ACQ_CORE_STA_FSM_STATE_OFFSET 0
`define ACQ_CORE_STA_FSM_STATE 32'h00000007
`define ACQ_CORE_STA_FSM_ACQ_DONE_OFFSET 3
`define ACQ_CORE_STA_FSM_ACQ_DONE 32'h00000008
`define ACQ_CORE_STA_RESERVED1_OFFSET 4
`define ACQ_CORE_STA_RESERVED1 32'h000000f0
`define ACQ_CORE_STA_FC_TRANS_DONE_OFFSET 8
`define ACQ_CORE_STA_FC_TRANS_DONE 32'h00000100
`define ACQ_CORE_STA_FC_FULL_OFFSET 9
`define ACQ_CORE_STA_FC_FULL 32'h00000200
`define ACQ_CORE_STA_RESERVED2_OFFSET 10
`define ACQ_CORE_STA_RESERVED2 32'h0000fc00
`define ACQ_CORE_STA_DDR3_TRANS_DONE_OFFSET 16
`define ACQ_CORE_STA_DDR3_TRANS_DONE 32'h00010000
`define ACQ_CORE_STA_RESERVED3_OFFSET 17
`define ACQ_CORE_STA_RESERVED3 32'hfffe0000
`define ADDR_ACQ_CORE_TRIG_CFG         8'h8
`define ACQ_CORE_TRIG_CFG_HW_TRIG_SEL_OFFSET 0
`define ACQ_CORE_TRIG_CFG_HW_TRIG_SEL 32'h00000001
`define ACQ_CORE_TRIG_CFG_HW_TRIG_POL_OFFSET 1
`define ACQ_CORE_TRIG_CFG_HW_TRIG_POL 32'h00000002
`define ACQ_CORE_TRIG_CFG_HW_TRIG_EN_OFFSET 2
`define ACQ_CORE_TRIG_CFG_HW_TRIG_EN 32'h00000004
`define ACQ_CORE_TRIG_CFG_SW_TRIG_EN_OFFSET 3
`define ACQ_CORE_TRIG_CFG_SW_TRIG_EN 32'h00000008
`define ACQ_CORE_TRIG_CFG_INT_TRIG_SEL_OFFSET 4
`define ACQ_CORE_TRIG_CFG_INT_TRIG_SEL 32'h000001f0
`define ACQ_CORE_TRIG_CFG_RESERVED_OFFSET 9
`define ACQ_CORE_TRIG_CFG_RESERVED 32'hfffffe00
`define ADDR_ACQ_CORE_TRIG_DATA_CFG    8'hc
`define ACQ_CORE_TRIG_DATA_CFG_THRES_FILT_OFFSET 0
`define ACQ_CORE_TRIG_DATA_CFG_THRES_FILT 32'h000000ff
`define ACQ_CORE_TRIG_DATA_CFG_RESERVED_OFFSET 8
`define ACQ_CORE_TRIG_DATA_CFG_RESERVED 32'hffffff00
`define ADDR_ACQ_CORE_TRIG_DATA_THRES  8'h10
`define ADDR_ACQ_CORE_TRIG_DLY         8'h14
`define ADDR_ACQ_CORE_SW_TRIG          8'h18
`define ADDR_ACQ_CORE_SHOTS            8'h1c
`define ACQ_CORE_SHOTS_NB_OFFSET 0
`define ACQ_CORE_SHOTS_NB 32'h0000ffff
`define ACQ_CORE_SHOTS_RESERVED_OFFSET 16
`define ACQ_CORE_SHOTS_RESERVED 32'hffff0000
`define ADDR_ACQ_CORE_TRIG_POS         8'h20
`define ADDR_ACQ_CORE_PRE_SAMPLES      8'h24
`define ADDR_ACQ_CORE_POST_SAMPLES     8'h28
`define ADDR_ACQ_CORE_SAMPLES_CNT      8'h2c
`define ADDR_ACQ_CORE_DDR3_START_ADDR  8'h30
`define ADDR_ACQ_CORE_DDR3_END_ADDR    8'h34
`define ADDR_ACQ_CORE_ACQ_CHAN_CTL     8'h38
`define ACQ_CORE_ACQ_CHAN_CTL_WHICH_OFFSET 0
`define ACQ_CORE_ACQ_CHAN_CTL_WHICH 32'h0000001f
`define ACQ_CORE_ACQ_CHAN_CTL_RESERVED_OFFSET 5
`define ACQ_CORE_ACQ_CHAN_CTL_RESERVED 32'h000000e0
`define ACQ_CORE_ACQ_CHAN_CTL_DTRIG_WHICH_OFFSET 8
`define ACQ_CORE_ACQ_CHAN_CTL_DTRIG_WHICH 32'h00001f00
`define ACQ_CORE_ACQ_CHAN_CTL_RESERVED1_OFFSET 13
`define ACQ_CORE_ACQ_CHAN_CTL_RESERVED1 32'hffffe000
`define ADDR_ACQ_CORE_CH0_DESC         8'h3c
`define ACQ_CORE_CH0_DESC_INT_WIDTH_OFFSET 0
`define ACQ_CORE_CH0_DESC_INT_WIDTH 32'h0000ffff
`define ACQ_CORE_CH0_DESC_NUM_COALESCE_OFFSET 16
`define ACQ_CORE_CH0_DESC_NUM_COALESCE 32'hffff0000
`define ADDR_ACQ_CORE_CH0_ATOM_DESC    8'h40
`define ACQ_CORE_CH0_ATOM_DESC_NUM_ATOMS_OFFSET 0
`define ACQ_CORE_CH0_ATOM_DESC_NUM_ATOMS 32'h0000ffff
`define ACQ_CORE_CH0_ATOM_DESC_ATOM_WIDTH_OFFSET 16
`define ACQ_CORE_CH0_ATOM_DESC_ATOM_WIDTH 32'hffff0000
`define ADDR_ACQ_CORE_CH1_DESC         8'h44
`define ACQ_CORE_CH1_DESC_INT_WIDTH_OFFSET 0
`define ACQ_CORE_CH1_DESC_INT_WIDTH 32'h0000ffff
`define ACQ_CORE_CH1_DESC_NUM_COALESCE_OFFSET 16
`define ACQ_CORE_CH1_DESC_NUM_COALESCE 32'hffff0000
`define ADDR_ACQ_CORE_CH1_ATOM_DESC    8'h48
`define ACQ_CORE_CH1_ATOM_DESC_NUM_ATOMS_OFFSET 0
`define ACQ_CORE_CH1_ATOM_DESC_NUM_ATOMS 32'h0000ffff
`define ACQ_CORE_CH1_ATOM_DESC_ATOM_WIDTH_OFFSET 16
`define ACQ_CORE_CH1_ATOM_DESC_ATOM_WIDTH 32'hffff0000
`define ADDR_ACQ_CORE_CH2_DESC         8'h4c
`define ACQ_CORE_CH2_DESC_INT_WIDTH_OFFSET 0
`define ACQ_CORE_CH2_DESC_INT_WIDTH 32'h0000ffff
`define ACQ_CORE_CH2_DESC_NUM_COALESCE_OFFSET 16
`define ACQ_CORE_CH2_DESC_NUM_COALESCE 32'hffff0000
`define ADDR_ACQ_CORE_CH2_ATOM_DESC    8'h50
`define ACQ_CORE_CH2_ATOM_DESC_NUM_ATOMS_OFFSET 0
`define ACQ_CORE_CH2_ATOM_DESC_NUM_ATOMS 32'h0000ffff
`define ACQ_CORE_CH2_ATOM_DESC_ATOM_WIDTH_OFFSET 16
`define ACQ_CORE_CH2_ATOM_DESC_ATOM_WIDTH 32'hffff0000
`define ADDR_ACQ_CORE_CH3_DESC         8'h54
`define ACQ_CORE_CH3_DESC_INT_WIDTH_OFFSET 0
`define ACQ_CORE_CH3_DESC_INT_WIDTH 32'h0000ffff
`define ACQ_CORE_CH3_DESC_NUM_COALESCE_OFFSET 16
`define ACQ_CORE_CH3_DESC_NUM_COALESCE 32'hffff0000
`define ADDR_ACQ_CORE_CH3_ATOM_DESC    8'h58
`define ACQ_CORE_CH3_ATOM_DESC_NUM_ATOMS_OFFSET 0
`define ACQ_CORE_CH3_ATOM_DESC_NUM_ATOMS 32'h0000ffff
`define ACQ_CORE_CH3_ATOM_DESC_ATOM_WIDTH_OFFSET 16
`define ACQ_CORE_CH3_ATOM_DESC_ATOM_WIDTH 32'hffff0000
`define ADDR_ACQ_CORE_CH4_DESC         8'h5c
`define ACQ_CORE_CH4_DESC_INT_WIDTH_OFFSET 0
`define ACQ_CORE_CH4_DESC_INT_WIDTH 32'h0000ffff
`define ACQ_CORE_CH4_DESC_NUM_COALESCE_OFFSET 16
`define ACQ_CORE_CH4_DESC_NUM_COALESCE 32'hffff0000
`define ADDR_ACQ_CORE_CH4_ATOM_DESC    8'h60
`define ACQ_CORE_CH4_ATOM_DESC_NUM_ATOMS_OFFSET 0
`define ACQ_CORE_CH4_ATOM_DESC_NUM_ATOMS 32'h0000ffff
`define ACQ_CORE_CH4_ATOM_DESC_ATOM_WIDTH_OFFSET 16
`define ACQ_CORE_CH4_ATOM_DESC_ATOM_WIDTH 32'hffff0000
`define ADDR_ACQ_CORE_CH5_DESC         8'h64
`define ACQ_CORE_CH5_DESC_INT_WIDTH_OFFSET 0
`define ACQ_CORE_CH5_DESC_INT_WIDTH 32'h0000ffff
`define ACQ_CORE_CH5_DESC_NUM_COALESCE_OFFSET 16
`define ACQ_CORE_CH5_DESC_NUM_COALESCE 32'hffff0000
`define ADDR_ACQ_CORE_CH5_ATOM_DESC    8'h68
`define ACQ_CORE_CH5_ATOM_DESC_NUM_ATOMS_OFFSET 0
`define ACQ_CORE_CH5_ATOM_DESC_NUM_ATOMS 32'h0000ffff
`define ACQ_CORE_CH5_ATOM_DESC_ATOM_WIDTH_OFFSET 16
`define ACQ_CORE_CH5_ATOM_DESC_ATOM_WIDTH 32'hffff0000
`define ADDR_ACQ_CORE_CH6_DESC         8'h6c
`define ACQ_CORE_CH6_DESC_INT_WIDTH_OFFSET 0
`define ACQ_CORE_CH6_DESC_INT_WIDTH 32'h0000ffff
`define ACQ_CORE_CH6_DESC_NUM_COALESCE_OFFSET 16
`define ACQ_CORE_CH6_DESC_NUM_COALESCE 32'hffff0000
`define ADDR_ACQ_CORE_CH6_ATOM_DESC    8'h70
`define ACQ_CORE_CH6_ATOM_DESC_NUM_ATOMS_OFFSET 0
`define ACQ_CORE_CH6_ATOM_DESC_NUM_ATOMS 32'h0000ffff
`define ACQ_CORE_CH6_ATOM_DESC_ATOM_WIDTH_OFFSET 16
`define ACQ_CORE_CH6_ATOM_DESC_ATOM_WIDTH 32'hffff0000
`define ADDR_ACQ_CORE_CH7_DESC         8'h74
`define ACQ_CORE_CH7_DESC_INT_WIDTH_OFFSET 0
`define ACQ_CORE_CH7_DESC_INT_WIDTH 32'h0000ffff
`define ACQ_CORE_CH7_DESC_NUM_COALESCE_OFFSET 16
`define ACQ_CORE_CH7_DESC_NUM_COALESCE 32'hffff0000
`define ADDR_ACQ_CORE_CH7_ATOM_DESC    8'h78
`define ACQ_CORE_CH7_ATOM_DESC_NUM_ATOMS_OFFSET 0
`define ACQ_CORE_CH7_ATOM_DESC_NUM_ATOMS 32'h0000ffff
`define ACQ_CORE_CH7_ATOM_DESC_ATOM_WIDTH_OFFSET 16
`define ACQ_CORE_CH7_ATOM_DESC_ATOM_WIDTH 32'hffff0000
`define ADDR_ACQ_CORE_CH8_DESC         8'h7c
`define ACQ_CORE_CH8_DESC_INT_WIDTH_OFFSET 0
`define ACQ_CORE_CH8_DESC_INT_WIDTH 32'h0000ffff
`define ACQ_CORE_CH8_DESC_NUM_COALESCE_OFFSET 16
`define ACQ_CORE_CH8_DESC_NUM_COALESCE 32'hffff0000
`define ADDR_ACQ_CORE_CH8_ATOM_DESC    8'h80
`define ACQ_CORE_CH8_ATOM_DESC_NUM_ATOMS_OFFSET 0
`define ACQ_CORE_CH8_ATOM_DESC_NUM_ATOMS 32'h0000ffff
`define ACQ_CORE_CH8_ATOM_DESC_ATOM_WIDTH_OFFSET 16
`define ACQ_CORE_CH8_ATOM_DESC_ATOM_WIDTH 32'hffff0000
`define ADDR_ACQ_CORE_CH9_DESC         8'h84
`define ACQ_CORE_CH9_DESC_INT_WIDTH_OFFSET 0
`define ACQ_CORE_CH9_DESC_INT_WIDTH 32'h0000ffff
`define ACQ_CORE_CH9_DESC_NUM_COALESCE_OFFSET 16
`define ACQ_CORE_CH9_DESC_NUM_COALESCE 32'hffff0000
`define ADDR_ACQ_CORE_CH9_ATOM_DESC    8'h88
`define ACQ_CORE_CH9_ATOM_DESC_NUM_ATOMS_OFFSET 0
`define ACQ_CORE_CH9_ATOM_DESC_NUM_ATOMS 32'h0000ffff
`define ACQ_CORE_CH9_ATOM_DESC_ATOM_WIDTH_OFFSET 16
`define ACQ_CORE_CH9_ATOM_DESC_ATOM_WIDTH 32'hffff0000
`define ADDR_ACQ_CORE_CH10_DESC        8'h8c
`define ACQ_CORE_CH10_DESC_INT_WIDTH_OFFSET 0
`define ACQ_CORE_CH10_DESC_INT_WIDTH 32'h0000ffff
`define ACQ_CORE_CH10_DESC_NUM_COALESCE_OFFSET 16
`define ACQ_CORE_CH10_DESC_NUM_COALESCE 32'hffff0000
`define ADDR_ACQ_CORE_CH10_ATOM_DESC   8'h90
`define ACQ_CORE_CH10_ATOM_DESC_NUM_ATOMS_OFFSET 0
`define ACQ_CORE_CH10_ATOM_DESC_NUM_ATOMS 32'h0000ffff
`define ACQ_CORE_CH10_ATOM_DESC_ATOM_WIDTH_OFFSET 16
`define ACQ_CORE_CH10_ATOM_DESC_ATOM_WIDTH 32'hffff0000
`define ADDR_ACQ_CORE_CH11_DESC        8'h94
`define ACQ_CORE_CH11_DESC_INT_WIDTH_OFFSET 0
`define ACQ_CORE_CH11_DESC_INT_WIDTH 32'h0000ffff
`define ACQ_CORE_CH11_DESC_NUM_COALESCE_OFFSET 16
`define ACQ_CORE_CH11_DESC_NUM_COALESCE 32'hffff0000
`define ADDR_ACQ_CORE_CH11_ATOM_DESC   8'h98
`define ACQ_CORE_CH11_ATOM_DESC_NUM_ATOMS_OFFSET 0
`define ACQ_CORE_CH11_ATOM_DESC_NUM_ATOMS 32'h0000ffff
`define ACQ_CORE_CH11_ATOM_DESC_ATOM_WIDTH_OFFSET 16
`define ACQ_CORE_CH11_ATOM_DESC_ATOM_WIDTH 32'hffff0000
`define ADDR_ACQ_CORE_CH12_DESC        8'h9c
`define ACQ_CORE_CH12_DESC_INT_WIDTH_OFFSET 0
`define ACQ_CORE_CH12_DESC_INT_WIDTH 32'h0000ffff
`define ACQ_CORE_CH12_DESC_NUM_COALESCE_OFFSET 16
`define ACQ_CORE_CH12_DESC_NUM_COALESCE 32'hffff0000
`define ADDR_ACQ_CORE_CH12_ATOM_DESC   8'ha0
`define ACQ_CORE_CH12_ATOM_DESC_NUM_ATOMS_OFFSET 0
`define ACQ_CORE_CH12_ATOM_DESC_NUM_ATOMS 32'h0000ffff
`define ACQ_CORE_CH12_ATOM_DESC_ATOM_WIDTH_OFFSET 16
`define ACQ_CORE_CH12_ATOM_DESC_ATOM_WIDTH 32'hffff0000
`define ADDR_ACQ_CORE_CH13_DESC        8'ha4
`define ACQ_CORE_CH13_DESC_INT_WIDTH_OFFSET 0
`define ACQ_CORE_CH13_DESC_INT_WIDTH 32'h0000ffff
`define ACQ_CORE_CH13_DESC_NUM_COALESCE_OFFSET 16
`define ACQ_CORE_CH13_DESC_NUM_COALESCE 32'hffff0000
`define ADDR_ACQ_CORE_CH13_ATOM_DESC   8'ha8
`define ACQ_CORE_CH13_ATOM_DESC_NUM_ATOMS_OFFSET 0
`define ACQ_CORE_CH13_ATOM_DESC_NUM_ATOMS 32'h0000ffff
`define ACQ_CORE_CH13_ATOM_DESC_ATOM_WIDTH_OFFSET 16
`define ACQ_CORE_CH13_ATOM_DESC_ATOM_WIDTH 32'hffff0000
`define ADDR_ACQ_CORE_CH14_DESC        8'hac
`define ACQ_CORE_CH14_DESC_INT_WIDTH_OFFSET 0
`define ACQ_CORE_CH14_DESC_INT_WIDTH 32'h0000ffff
`define ACQ_CORE_CH14_DESC_NUM_COALESCE_OFFSET 16
`define ACQ_CORE_CH14_DESC_NUM_COALESCE 32'hffff0000
`define ADDR_ACQ_CORE_CH14_ATOM_DESC   8'hb0
`define ACQ_CORE_CH14_ATOM_DESC_NUM_ATOMS_OFFSET 0
`define ACQ_CORE_CH14_ATOM_DESC_NUM_ATOMS 32'h0000ffff
`define ACQ_CORE_CH14_ATOM_DESC_ATOM_WIDTH_OFFSET 16
`define ACQ_CORE_CH14_ATOM_DESC_ATOM_WIDTH 32'hffff0000
`define ADDR_ACQ_CORE_CH15_DESC        8'hb4
`define ACQ_CORE_CH15_DESC_INT_WIDTH_OFFSET 0
`define ACQ_CORE_CH15_DESC_INT_WIDTH 32'h0000ffff
`define ACQ_CORE_CH15_DESC_NUM_COALESCE_OFFSET 16
`define ACQ_CORE_CH15_DESC_NUM_COALESCE 32'hffff0000
`define ADDR_ACQ_CORE_CH15_ATOM_DESC   8'hb8
`define ACQ_CORE_CH15_ATOM_DESC_NUM_ATOMS_OFFSET 0
`define ACQ_CORE_CH15_ATOM_DESC_NUM_ATOMS 32'h0000ffff
`define ACQ_CORE_CH15_ATOM_DESC_ATOM_WIDTH_OFFSET 16
`define ACQ_CORE_CH15_ATOM_DESC_ATOM_WIDTH 32'hffff0000
`define ADDR_ACQ_CORE_CH16_DESC        8'hbc
`define ACQ_CORE_CH16_DESC_INT_WIDTH_OFFSET 0
`define ACQ_CORE_CH16_DESC_INT_WIDTH 32'h0000ffff
`define ACQ_CORE_CH16_DESC_NUM_COALESCE_OFFSET 16
`define ACQ_CORE_CH16_DESC_NUM_COALESCE 32'hffff0000
`define ADDR_ACQ_CORE_CH16_ATOM_DESC   8'hc0
`define ACQ_CORE_CH16_ATOM_DESC_NUM_ATOMS_OFFSET 0
`define ACQ_CORE_CH16_ATOM_DESC_NUM_ATOMS 32'h0000ffff
`define ACQ_CORE_CH16_ATOM_DESC_ATOM_WIDTH_OFFSET 16
`define ACQ_CORE_CH16_ATOM_DESC_ATOM_WIDTH 32'hffff0000
`define ADDR_ACQ_CORE_CH17_DESC        8'hc4
`define ACQ_CORE_CH17_DESC_INT_WIDTH_OFFSET 0
`define ACQ_CORE_CH17_DESC_INT_WIDTH 32'h0000ffff
`define ACQ_CORE_CH17_DESC_NUM_COALESCE_OFFSET 16
`define ACQ_CORE_CH17_DESC_NUM_COALESCE 32'hffff0000
`define ADDR_ACQ_CORE_CH17_ATOM_DESC   8'hc8
`define ACQ_CORE_CH17_ATOM_DESC_NUM_ATOMS_OFFSET 0
`define ACQ_CORE_CH17_ATOM_DESC_NUM_ATOMS 32'h0000ffff
`define ACQ_CORE_CH17_ATOM_DESC_ATOM_WIDTH_OFFSET 16
`define ACQ_CORE_CH17_ATOM_DESC_ATOM_WIDTH 32'hffff0000
`define ADDR_ACQ_CORE_CH18_DESC        8'hcc
`define ACQ_CORE_CH18_DESC_INT_WIDTH_OFFSET 0
`define ACQ_CORE_CH18_DESC_INT_WIDTH 32'h0000ffff
`define ACQ_CORE_CH18_DESC_NUM_COALESCE_OFFSET 16
`define ACQ_CORE_CH18_DESC_NUM_COALESCE 32'hffff0000
`define ADDR_ACQ_CORE_CH18_ATOM_DESC   8'hd0
`define ACQ_CORE_CH18_ATOM_DESC_NUM_ATOMS_OFFSET 0
`define ACQ_CORE_CH18_ATOM_DESC_NUM_ATOMS 32'h0000ffff
`define ACQ_CORE_CH18_ATOM_DESC_ATOM_WIDTH_OFFSET 16
`define ACQ_CORE_CH18_ATOM_DESC_ATOM_WIDTH 32'hffff0000
`define ADDR_ACQ_CORE_CH19_DESC        8'hd4
`define ACQ_CORE_CH19_DESC_INT_WIDTH_OFFSET 0
`define ACQ_CORE_CH19_DESC_INT_WIDTH 32'h0000ffff
`define ACQ_CORE_CH19_DESC_NUM_COALESCE_OFFSET 16
`define ACQ_CORE_CH19_DESC_NUM_COALESCE 32'hffff0000
`define ADDR_ACQ_CORE_CH19_ATOM_DESC   8'hd8
`define ACQ_CORE_CH19_ATOM_DESC_NUM_ATOMS_OFFSET 0
`define ACQ_CORE_CH19_ATOM_DESC_NUM_ATOMS 32'h0000ffff
`define ACQ_CORE_CH19_ATOM_DESC_ATOM_WIDTH_OFFSET 16
`define ACQ_CORE_CH19_ATOM_DESC_ATOM_WIDTH 32'hffff0000
`define ADDR_ACQ_CORE_CH20_DESC        8'hdc
`define ACQ_CORE_CH20_DESC_INT_WIDTH_OFFSET 0
`define ACQ_CORE_CH20_DESC_INT_WIDTH 32'h0000ffff
`define ACQ_CORE_CH20_DESC_NUM_COALESCE_OFFSET 16
`define ACQ_CORE_CH20_DESC_NUM_COALESCE 32'hffff0000
`define ADDR_ACQ_CORE_CH20_ATOM_DESC   8'he0
`define ACQ_CORE_CH20_ATOM_DESC_NUM_ATOMS_OFFSET 0
`define ACQ_CORE_CH20_ATOM_DESC_NUM_ATOMS 32'h0000ffff
`define ACQ_CORE_CH20_ATOM_DESC_ATOM_WIDTH_OFFSET 16
`define ACQ_CORE_CH20_ATOM_DESC_ATOM_WIDTH 32'hffff0000
`define ADDR_ACQ_CORE_CH21_DESC        8'he4
`define ACQ_CORE_CH21_DESC_INT_WIDTH_OFFSET 0
`define ACQ_CORE_CH21_DESC_INT_WIDTH 32'h0000ffff
`define ACQ_CORE_CH21_DESC_NUM_COALESCE_OFFSET 16
`define ACQ_CORE_CH21_DESC_NUM_COALESCE 32'hffff0000
`define ADDR_ACQ_CORE_CH21_ATOM_DESC   8'he8
`define ACQ_CORE_CH21_ATOM_DESC_NUM_ATOMS_OFFSET 0
`define ACQ_CORE_CH21_ATOM_DESC_NUM_ATOMS 32'h0000ffff
`define ACQ_CORE_CH21_ATOM_DESC_ATOM_WIDTH_OFFSET 16
`define ACQ_CORE_CH21_ATOM_DESC_ATOM_WIDTH 32'hffff0000
`define ADDR_ACQ_CORE_CH22_DESC        8'hec
`define ACQ_CORE_CH22_DESC_INT_WIDTH_OFFSET 0
`define ACQ_CORE_CH22_DESC_INT_WIDTH 32'h0000ffff
`define ACQ_CORE_CH22_DESC_NUM_COALESCE_OFFSET 16
`define ACQ_CORE_CH22_DESC_NUM_COALESCE 32'hffff0000
`define ADDR_ACQ_CORE_CH22_ATOM_DESC   8'hf0
`define ACQ_CORE_CH22_ATOM_DESC_NUM_ATOMS_OFFSET 0
`define ACQ_CORE_CH22_ATOM_DESC_NUM_ATOMS 32'h0000ffff
`define ACQ_CORE_CH22_ATOM_DESC_ATOM_WIDTH_OFFSET 16
`define ACQ_CORE_CH22_ATOM_DESC_ATOM_WIDTH 32'hffff0000
`define ADDR_ACQ_CORE_CH23_DESC        8'hf4
`define ACQ_CORE_CH23_DESC_INT_WIDTH_OFFSET 0
`define ACQ_CORE_CH23_DESC_INT_WIDTH 32'h0000ffff
`define ACQ_CORE_CH23_DESC_NUM_COALESCE_OFFSET 16
`define ACQ_CORE_CH23_DESC_NUM_COALESCE 32'hffff0000
`define ADDR_ACQ_CORE_CH23_ATOM_DESC   8'hf8
`define ACQ_CORE_CH23_ATOM_DESC_NUM_ATOMS_OFFSET 0
`define ACQ_CORE_CH23_ATOM_DESC_NUM_ATOMS 32'h0000ffff
`define ACQ_CORE_CH23_ATOM_DESC_ATOM_WIDTH_OFFSET 16
`define ACQ_CORE_CH23_ATOM_DESC_ATOM_WIDTH 32'hffff0000
