`define ADDR_WB_FMC_ADC_COMMON_CSR_FMC_STATUS 4'h0
`define WB_FMC_ADC_COMMON_CSR_FMC_STATUS_MMCM_LOCKED_OFFSET 0
`define WB_FMC_ADC_COMMON_CSR_FMC_STATUS_MMCM_LOCKED 32'h00000001
`define WB_FMC_ADC_COMMON_CSR_FMC_STATUS_PWR_GOOD_OFFSET 1
`define WB_FMC_ADC_COMMON_CSR_FMC_STATUS_PWR_GOOD 32'h00000002
`define WB_FMC_ADC_COMMON_CSR_FMC_STATUS_PRST_OFFSET 2
`define WB_FMC_ADC_COMMON_CSR_FMC_STATUS_PRST 32'h00000004
`define WB_FMC_ADC_COMMON_CSR_FMC_STATUS_RESERVED_OFFSET 3
`define WB_FMC_ADC_COMMON_CSR_FMC_STATUS_RESERVED 32'h7ffffff8
`define ADDR_WB_FMC_ADC_COMMON_CSR_TRIGGER 4'h4
`define WB_FMC_ADC_COMMON_CSR_TRIGGER_DIR_OFFSET 0
`define WB_FMC_ADC_COMMON_CSR_TRIGGER_DIR 32'h00000001
`define WB_FMC_ADC_COMMON_CSR_TRIGGER_TERM_OFFSET 1
`define WB_FMC_ADC_COMMON_CSR_TRIGGER_TERM 32'h00000002
`define WB_FMC_ADC_COMMON_CSR_TRIGGER_TRIG_VAL_OFFSET 2
`define WB_FMC_ADC_COMMON_CSR_TRIGGER_TRIG_VAL 32'h00000004
`define WB_FMC_ADC_COMMON_CSR_TRIGGER_RESERVED_OFFSET 3
`define WB_FMC_ADC_COMMON_CSR_TRIGGER_RESERVED 32'hfffffff8
`define ADDR_WB_FMC_ADC_COMMON_CSR_MONITOR 4'h8
`define WB_FMC_ADC_COMMON_CSR_MONITOR_TEST_DATA_EN_OFFSET 0
`define WB_FMC_ADC_COMMON_CSR_MONITOR_TEST_DATA_EN 32'h00000001
`define WB_FMC_ADC_COMMON_CSR_MONITOR_LED1_OFFSET 1
`define WB_FMC_ADC_COMMON_CSR_MONITOR_LED1 32'h00000002
`define WB_FMC_ADC_COMMON_CSR_MONITOR_LED2_OFFSET 2
`define WB_FMC_ADC_COMMON_CSR_MONITOR_LED2 32'h00000004
`define WB_FMC_ADC_COMMON_CSR_MONITOR_LED3_OFFSET 3
`define WB_FMC_ADC_COMMON_CSR_MONITOR_LED3 32'h00000008
`define WB_FMC_ADC_COMMON_CSR_MONITOR_MMCM_RST_OFFSET 4
`define WB_FMC_ADC_COMMON_CSR_MONITOR_MMCM_RST 32'h00000010
`define WB_FMC_ADC_COMMON_CSR_MONITOR_RESERVED_OFFSET 5
`define WB_FMC_ADC_COMMON_CSR_MONITOR_RESERVED 32'hffffffe0
