`define ADDR_WB_TRIG_MUX_CH0_CTL       8'h0
`define WB_TRIG_MUX_CH0_CTL_RCV_SRC_OFFSET 0
`define WB_TRIG_MUX_CH0_CTL_RCV_SRC 32'h00000001
`define WB_TRIG_MUX_CH0_CTL_RCV_IN_SEL_OFFSET 8
`define WB_TRIG_MUX_CH0_CTL_RCV_IN_SEL 32'h0000ff00
`define WB_TRIG_MUX_CH0_CTL_TRANSM_SRC_OFFSET 16
`define WB_TRIG_MUX_CH0_CTL_TRANSM_SRC 32'h00010000
`define WB_TRIG_MUX_CH0_CTL_TRANSM_OUT_SEL_OFFSET 24
`define WB_TRIG_MUX_CH0_CTL_TRANSM_OUT_SEL 32'hff000000
`define ADDR_WB_TRIG_MUX_CH0_DUMMY     8'h4
`define ADDR_WB_TRIG_MUX_CH1_CTL       8'h8
`define WB_TRIG_MUX_CH1_CTL_RCV_SRC_OFFSET 0
`define WB_TRIG_MUX_CH1_CTL_RCV_SRC 32'h00000001
`define WB_TRIG_MUX_CH1_CTL_RCV_IN_SEL_OFFSET 8
`define WB_TRIG_MUX_CH1_CTL_RCV_IN_SEL 32'h0000ff00
`define WB_TRIG_MUX_CH1_CTL_TRANSM_SRC_OFFSET 16
`define WB_TRIG_MUX_CH1_CTL_TRANSM_SRC 32'h00010000
`define WB_TRIG_MUX_CH1_CTL_TRANSM_OUT_SEL_OFFSET 24
`define WB_TRIG_MUX_CH1_CTL_TRANSM_OUT_SEL 32'hff000000
`define ADDR_WB_TRIG_MUX_CH1_DUMMY     8'hc
`define ADDR_WB_TRIG_MUX_CH2_CTL       8'h10
`define WB_TRIG_MUX_CH2_CTL_RCV_SRC_OFFSET 0
`define WB_TRIG_MUX_CH2_CTL_RCV_SRC 32'h00000001
`define WB_TRIG_MUX_CH2_CTL_RCV_IN_SEL_OFFSET 8
`define WB_TRIG_MUX_CH2_CTL_RCV_IN_SEL 32'h0000ff00
`define WB_TRIG_MUX_CH2_CTL_TRANSM_SRC_OFFSET 16
`define WB_TRIG_MUX_CH2_CTL_TRANSM_SRC 32'h00010000
`define WB_TRIG_MUX_CH2_CTL_TRANSM_OUT_SEL_OFFSET 24
`define WB_TRIG_MUX_CH2_CTL_TRANSM_OUT_SEL 32'hff000000
`define ADDR_WB_TRIG_MUX_CH2_DUMMY     8'h14
`define ADDR_WB_TRIG_MUX_CH3_CTL       8'h18
`define WB_TRIG_MUX_CH3_CTL_RCV_SRC_OFFSET 0
`define WB_TRIG_MUX_CH3_CTL_RCV_SRC 32'h00000001
`define WB_TRIG_MUX_CH3_CTL_RCV_IN_SEL_OFFSET 8
`define WB_TRIG_MUX_CH3_CTL_RCV_IN_SEL 32'h0000ff00
`define WB_TRIG_MUX_CH3_CTL_TRANSM_SRC_OFFSET 16
`define WB_TRIG_MUX_CH3_CTL_TRANSM_SRC 32'h00010000
`define WB_TRIG_MUX_CH3_CTL_TRANSM_OUT_SEL_OFFSET 24
`define WB_TRIG_MUX_CH3_CTL_TRANSM_OUT_SEL 32'hff000000
`define ADDR_WB_TRIG_MUX_CH3_DUMMY     8'h1c
`define ADDR_WB_TRIG_MUX_CH4_CTL       8'h20
`define WB_TRIG_MUX_CH4_CTL_RCV_SRC_OFFSET 0
`define WB_TRIG_MUX_CH4_CTL_RCV_SRC 32'h00000001
`define WB_TRIG_MUX_CH4_CTL_RCV_IN_SEL_OFFSET 8
`define WB_TRIG_MUX_CH4_CTL_RCV_IN_SEL 32'h0000ff00
`define WB_TRIG_MUX_CH4_CTL_TRANSM_SRC_OFFSET 16
`define WB_TRIG_MUX_CH4_CTL_TRANSM_SRC 32'h00010000
`define WB_TRIG_MUX_CH4_CTL_TRANSM_OUT_SEL_OFFSET 24
`define WB_TRIG_MUX_CH4_CTL_TRANSM_OUT_SEL 32'hff000000
`define ADDR_WB_TRIG_MUX_CH4_DUMMY     8'h24
`define ADDR_WB_TRIG_MUX_CH5_CTL       8'h28
`define WB_TRIG_MUX_CH5_CTL_RCV_SRC_OFFSET 0
`define WB_TRIG_MUX_CH5_CTL_RCV_SRC 32'h00000001
`define WB_TRIG_MUX_CH5_CTL_RCV_IN_SEL_OFFSET 8
`define WB_TRIG_MUX_CH5_CTL_RCV_IN_SEL 32'h0000ff00
`define WB_TRIG_MUX_CH5_CTL_TRANSM_SRC_OFFSET 16
`define WB_TRIG_MUX_CH5_CTL_TRANSM_SRC 32'h00010000
`define WB_TRIG_MUX_CH5_CTL_TRANSM_OUT_SEL_OFFSET 24
`define WB_TRIG_MUX_CH5_CTL_TRANSM_OUT_SEL 32'hff000000
`define ADDR_WB_TRIG_MUX_CH5_DUMMY     8'h2c
`define ADDR_WB_TRIG_MUX_CH6_CTL       8'h30
`define WB_TRIG_MUX_CH6_CTL_RCV_SRC_OFFSET 0
`define WB_TRIG_MUX_CH6_CTL_RCV_SRC 32'h00000001
`define WB_TRIG_MUX_CH6_CTL_RCV_IN_SEL_OFFSET 8
`define WB_TRIG_MUX_CH6_CTL_RCV_IN_SEL 32'h0000ff00
`define WB_TRIG_MUX_CH6_CTL_TRANSM_SRC_OFFSET 16
`define WB_TRIG_MUX_CH6_CTL_TRANSM_SRC 32'h00010000
`define WB_TRIG_MUX_CH6_CTL_TRANSM_OUT_SEL_OFFSET 24
`define WB_TRIG_MUX_CH6_CTL_TRANSM_OUT_SEL 32'hff000000
`define ADDR_WB_TRIG_MUX_CH6_DUMMY     8'h34
`define ADDR_WB_TRIG_MUX_CH7_CTL       8'h38
`define WB_TRIG_MUX_CH7_CTL_RCV_SRC_OFFSET 0
`define WB_TRIG_MUX_CH7_CTL_RCV_SRC 32'h00000001
`define WB_TRIG_MUX_CH7_CTL_RCV_IN_SEL_OFFSET 8
`define WB_TRIG_MUX_CH7_CTL_RCV_IN_SEL 32'h0000ff00
`define WB_TRIG_MUX_CH7_CTL_TRANSM_SRC_OFFSET 16
`define WB_TRIG_MUX_CH7_CTL_TRANSM_SRC 32'h00010000
`define WB_TRIG_MUX_CH7_CTL_TRANSM_OUT_SEL_OFFSET 24
`define WB_TRIG_MUX_CH7_CTL_TRANSM_OUT_SEL 32'hff000000
`define ADDR_WB_TRIG_MUX_CH7_DUMMY     8'h3c
`define ADDR_WB_TRIG_MUX_CH8_CTL       8'h40
`define WB_TRIG_MUX_CH8_CTL_RCV_SRC_OFFSET 0
`define WB_TRIG_MUX_CH8_CTL_RCV_SRC 32'h00000001
`define WB_TRIG_MUX_CH8_CTL_RCV_IN_SEL_OFFSET 8
`define WB_TRIG_MUX_CH8_CTL_RCV_IN_SEL 32'h0000ff00
`define WB_TRIG_MUX_CH8_CTL_TRANSM_SRC_OFFSET 16
`define WB_TRIG_MUX_CH8_CTL_TRANSM_SRC 32'h00010000
`define WB_TRIG_MUX_CH8_CTL_TRANSM_OUT_SEL_OFFSET 24
`define WB_TRIG_MUX_CH8_CTL_TRANSM_OUT_SEL 32'hff000000
`define ADDR_WB_TRIG_MUX_CH8_DUMMY     8'h44
`define ADDR_WB_TRIG_MUX_CH9_CTL       8'h48
`define WB_TRIG_MUX_CH9_CTL_RCV_SRC_OFFSET 0
`define WB_TRIG_MUX_CH9_CTL_RCV_SRC 32'h00000001
`define WB_TRIG_MUX_CH9_CTL_RCV_IN_SEL_OFFSET 8
`define WB_TRIG_MUX_CH9_CTL_RCV_IN_SEL 32'h0000ff00
`define WB_TRIG_MUX_CH9_CTL_TRANSM_SRC_OFFSET 16
`define WB_TRIG_MUX_CH9_CTL_TRANSM_SRC 32'h00010000
`define WB_TRIG_MUX_CH9_CTL_TRANSM_OUT_SEL_OFFSET 24
`define WB_TRIG_MUX_CH9_CTL_TRANSM_OUT_SEL 32'hff000000
`define ADDR_WB_TRIG_MUX_CH9_DUMMY     8'h4c
`define ADDR_WB_TRIG_MUX_CH10_CTL      8'h50
`define WB_TRIG_MUX_CH10_CTL_RCV_SRC_OFFSET 0
`define WB_TRIG_MUX_CH10_CTL_RCV_SRC 32'h00000001
`define WB_TRIG_MUX_CH10_CTL_RCV_IN_SEL_OFFSET 8
`define WB_TRIG_MUX_CH10_CTL_RCV_IN_SEL 32'h0000ff00
`define WB_TRIG_MUX_CH10_CTL_TRANSM_SRC_OFFSET 16
`define WB_TRIG_MUX_CH10_CTL_TRANSM_SRC 32'h00010000
`define WB_TRIG_MUX_CH10_CTL_TRANSM_OUT_SEL_OFFSET 24
`define WB_TRIG_MUX_CH10_CTL_TRANSM_OUT_SEL 32'hff000000
`define ADDR_WB_TRIG_MUX_CH10_DUMMY    8'h54
`define ADDR_WB_TRIG_MUX_CH11_CTL      8'h58
`define WB_TRIG_MUX_CH11_CTL_RCV_SRC_OFFSET 0
`define WB_TRIG_MUX_CH11_CTL_RCV_SRC 32'h00000001
`define WB_TRIG_MUX_CH11_CTL_RCV_IN_SEL_OFFSET 8
`define WB_TRIG_MUX_CH11_CTL_RCV_IN_SEL 32'h0000ff00
`define WB_TRIG_MUX_CH11_CTL_TRANSM_SRC_OFFSET 16
`define WB_TRIG_MUX_CH11_CTL_TRANSM_SRC 32'h00010000
`define WB_TRIG_MUX_CH11_CTL_TRANSM_OUT_SEL_OFFSET 24
`define WB_TRIG_MUX_CH11_CTL_TRANSM_OUT_SEL 32'hff000000
`define ADDR_WB_TRIG_MUX_CH11_DUMMY    8'h5c
`define ADDR_WB_TRIG_MUX_CH12_CTL      8'h60
`define WB_TRIG_MUX_CH12_CTL_RCV_SRC_OFFSET 0
`define WB_TRIG_MUX_CH12_CTL_RCV_SRC 32'h00000001
`define WB_TRIG_MUX_CH12_CTL_RCV_IN_SEL_OFFSET 8
`define WB_TRIG_MUX_CH12_CTL_RCV_IN_SEL 32'h0000ff00
`define WB_TRIG_MUX_CH12_CTL_TRANSM_SRC_OFFSET 16
`define WB_TRIG_MUX_CH12_CTL_TRANSM_SRC 32'h00010000
`define WB_TRIG_MUX_CH12_CTL_TRANSM_OUT_SEL_OFFSET 24
`define WB_TRIG_MUX_CH12_CTL_TRANSM_OUT_SEL 32'hff000000
`define ADDR_WB_TRIG_MUX_CH12_DUMMY    8'h64
`define ADDR_WB_TRIG_MUX_CH13_CTL      8'h68
`define WB_TRIG_MUX_CH13_CTL_RCV_SRC_OFFSET 0
`define WB_TRIG_MUX_CH13_CTL_RCV_SRC 32'h00000001
`define WB_TRIG_MUX_CH13_CTL_RCV_IN_SEL_OFFSET 8
`define WB_TRIG_MUX_CH13_CTL_RCV_IN_SEL 32'h0000ff00
`define WB_TRIG_MUX_CH13_CTL_TRANSM_SRC_OFFSET 16
`define WB_TRIG_MUX_CH13_CTL_TRANSM_SRC 32'h00010000
`define WB_TRIG_MUX_CH13_CTL_TRANSM_OUT_SEL_OFFSET 24
`define WB_TRIG_MUX_CH13_CTL_TRANSM_OUT_SEL 32'hff000000
`define ADDR_WB_TRIG_MUX_CH13_DUMMY    8'h6c
`define ADDR_WB_TRIG_MUX_CH14_CTL      8'h70
`define WB_TRIG_MUX_CH14_CTL_RCV_SRC_OFFSET 0
`define WB_TRIG_MUX_CH14_CTL_RCV_SRC 32'h00000001
`define WB_TRIG_MUX_CH14_CTL_RCV_IN_SEL_OFFSET 8
`define WB_TRIG_MUX_CH14_CTL_RCV_IN_SEL 32'h0000ff00
`define WB_TRIG_MUX_CH14_CTL_TRANSM_SRC_OFFSET 16
`define WB_TRIG_MUX_CH14_CTL_TRANSM_SRC 32'h00010000
`define WB_TRIG_MUX_CH14_CTL_TRANSM_OUT_SEL_OFFSET 24
`define WB_TRIG_MUX_CH14_CTL_TRANSM_OUT_SEL 32'hff000000
`define ADDR_WB_TRIG_MUX_CH14_DUMMY    8'h74
`define ADDR_WB_TRIG_MUX_CH15_CTL      8'h78
`define WB_TRIG_MUX_CH15_CTL_RCV_SRC_OFFSET 0
`define WB_TRIG_MUX_CH15_CTL_RCV_SRC 32'h00000001
`define WB_TRIG_MUX_CH15_CTL_RCV_IN_SEL_OFFSET 8
`define WB_TRIG_MUX_CH15_CTL_RCV_IN_SEL 32'h0000ff00
`define WB_TRIG_MUX_CH15_CTL_TRANSM_SRC_OFFSET 16
`define WB_TRIG_MUX_CH15_CTL_TRANSM_SRC 32'h00010000
`define WB_TRIG_MUX_CH15_CTL_TRANSM_OUT_SEL_OFFSET 24
`define WB_TRIG_MUX_CH15_CTL_TRANSM_OUT_SEL 32'hff000000
`define ADDR_WB_TRIG_MUX_CH15_DUMMY    8'h7c
`define ADDR_WB_TRIG_MUX_CH16_CTL      8'h80
`define WB_TRIG_MUX_CH16_CTL_RCV_SRC_OFFSET 0
`define WB_TRIG_MUX_CH16_CTL_RCV_SRC 32'h00000001
`define WB_TRIG_MUX_CH16_CTL_RCV_IN_SEL_OFFSET 8
`define WB_TRIG_MUX_CH16_CTL_RCV_IN_SEL 32'h0000ff00
`define WB_TRIG_MUX_CH16_CTL_TRANSM_SRC_OFFSET 16
`define WB_TRIG_MUX_CH16_CTL_TRANSM_SRC 32'h00010000
`define WB_TRIG_MUX_CH16_CTL_TRANSM_OUT_SEL_OFFSET 24
`define WB_TRIG_MUX_CH16_CTL_TRANSM_OUT_SEL 32'hff000000
`define ADDR_WB_TRIG_MUX_CH16_DUMMY    8'h84
`define ADDR_WB_TRIG_MUX_CH17_CTL      8'h88
`define WB_TRIG_MUX_CH17_CTL_RCV_SRC_OFFSET 0
`define WB_TRIG_MUX_CH17_CTL_RCV_SRC 32'h00000001
`define WB_TRIG_MUX_CH17_CTL_RCV_IN_SEL_OFFSET 8
`define WB_TRIG_MUX_CH17_CTL_RCV_IN_SEL 32'h0000ff00
`define WB_TRIG_MUX_CH17_CTL_TRANSM_SRC_OFFSET 16
`define WB_TRIG_MUX_CH17_CTL_TRANSM_SRC 32'h00010000
`define WB_TRIG_MUX_CH17_CTL_TRANSM_OUT_SEL_OFFSET 24
`define WB_TRIG_MUX_CH17_CTL_TRANSM_OUT_SEL 32'hff000000
`define ADDR_WB_TRIG_MUX_CH17_DUMMY    8'h8c
`define ADDR_WB_TRIG_MUX_CH18_CTL      8'h90
`define WB_TRIG_MUX_CH18_CTL_RCV_SRC_OFFSET 0
`define WB_TRIG_MUX_CH18_CTL_RCV_SRC 32'h00000001
`define WB_TRIG_MUX_CH18_CTL_RCV_IN_SEL_OFFSET 8
`define WB_TRIG_MUX_CH18_CTL_RCV_IN_SEL 32'h0000ff00
`define WB_TRIG_MUX_CH18_CTL_TRANSM_SRC_OFFSET 16
`define WB_TRIG_MUX_CH18_CTL_TRANSM_SRC 32'h00010000
`define WB_TRIG_MUX_CH18_CTL_TRANSM_OUT_SEL_OFFSET 24
`define WB_TRIG_MUX_CH18_CTL_TRANSM_OUT_SEL 32'hff000000
`define ADDR_WB_TRIG_MUX_CH18_DUMMY    8'h94
`define ADDR_WB_TRIG_MUX_CH19_CTL      8'h98
`define WB_TRIG_MUX_CH19_CTL_RCV_SRC_OFFSET 0
`define WB_TRIG_MUX_CH19_CTL_RCV_SRC 32'h00000001
`define WB_TRIG_MUX_CH19_CTL_RCV_IN_SEL_OFFSET 8
`define WB_TRIG_MUX_CH19_CTL_RCV_IN_SEL 32'h0000ff00
`define WB_TRIG_MUX_CH19_CTL_TRANSM_SRC_OFFSET 16
`define WB_TRIG_MUX_CH19_CTL_TRANSM_SRC 32'h00010000
`define WB_TRIG_MUX_CH19_CTL_TRANSM_OUT_SEL_OFFSET 24
`define WB_TRIG_MUX_CH19_CTL_TRANSM_OUT_SEL 32'hff000000
`define ADDR_WB_TRIG_MUX_CH19_DUMMY    8'h9c
`define ADDR_WB_TRIG_MUX_CH20_CTL      8'ha0
`define WB_TRIG_MUX_CH20_CTL_RCV_SRC_OFFSET 0
`define WB_TRIG_MUX_CH20_CTL_RCV_SRC 32'h00000001
`define WB_TRIG_MUX_CH20_CTL_RCV_IN_SEL_OFFSET 8
`define WB_TRIG_MUX_CH20_CTL_RCV_IN_SEL 32'h0000ff00
`define WB_TRIG_MUX_CH20_CTL_TRANSM_SRC_OFFSET 16
`define WB_TRIG_MUX_CH20_CTL_TRANSM_SRC 32'h00010000
`define WB_TRIG_MUX_CH20_CTL_TRANSM_OUT_SEL_OFFSET 24
`define WB_TRIG_MUX_CH20_CTL_TRANSM_OUT_SEL 32'hff000000
`define ADDR_WB_TRIG_MUX_CH20_DUMMY    8'ha4
`define ADDR_WB_TRIG_MUX_CH21_CTL      8'ha8
`define WB_TRIG_MUX_CH21_CTL_RCV_SRC_OFFSET 0
`define WB_TRIG_MUX_CH21_CTL_RCV_SRC 32'h00000001
`define WB_TRIG_MUX_CH21_CTL_RCV_IN_SEL_OFFSET 8
`define WB_TRIG_MUX_CH21_CTL_RCV_IN_SEL 32'h0000ff00
`define WB_TRIG_MUX_CH21_CTL_TRANSM_SRC_OFFSET 16
`define WB_TRIG_MUX_CH21_CTL_TRANSM_SRC 32'h00010000
`define WB_TRIG_MUX_CH21_CTL_TRANSM_OUT_SEL_OFFSET 24
`define WB_TRIG_MUX_CH21_CTL_TRANSM_OUT_SEL 32'hff000000
`define ADDR_WB_TRIG_MUX_CH21_DUMMY    8'hac
`define ADDR_WB_TRIG_MUX_CH22_CTL      8'hb0
`define WB_TRIG_MUX_CH22_CTL_RCV_SRC_OFFSET 0
`define WB_TRIG_MUX_CH22_CTL_RCV_SRC 32'h00000001
`define WB_TRIG_MUX_CH22_CTL_RCV_IN_SEL_OFFSET 8
`define WB_TRIG_MUX_CH22_CTL_RCV_IN_SEL 32'h0000ff00
`define WB_TRIG_MUX_CH22_CTL_TRANSM_SRC_OFFSET 16
`define WB_TRIG_MUX_CH22_CTL_TRANSM_SRC 32'h00010000
`define WB_TRIG_MUX_CH22_CTL_TRANSM_OUT_SEL_OFFSET 24
`define WB_TRIG_MUX_CH22_CTL_TRANSM_OUT_SEL 32'hff000000
`define ADDR_WB_TRIG_MUX_CH22_DUMMY    8'hb4
`define ADDR_WB_TRIG_MUX_CH23_CTL      8'hb8
`define WB_TRIG_MUX_CH23_CTL_RCV_SRC_OFFSET 0
`define WB_TRIG_MUX_CH23_CTL_RCV_SRC 32'h00000001
`define WB_TRIG_MUX_CH23_CTL_RCV_IN_SEL_OFFSET 8
`define WB_TRIG_MUX_CH23_CTL_RCV_IN_SEL 32'h0000ff00
`define WB_TRIG_MUX_CH23_CTL_TRANSM_SRC_OFFSET 16
`define WB_TRIG_MUX_CH23_CTL_TRANSM_SRC 32'h00010000
`define WB_TRIG_MUX_CH23_CTL_TRANSM_OUT_SEL_OFFSET 24
`define WB_TRIG_MUX_CH23_CTL_TRANSM_OUT_SEL 32'hff000000
`define ADDR_WB_TRIG_MUX_CH23_DUMMY    8'hbc
