`include "sample_tests1.vh"
`include "tf64_pcie_axi.vh"
