`define ADDR_WB_FMC_250M_4CH_CSR_FMC_STA 7'h0
`define WB_FMC_250M_4CH_CSR_FMC_STA_MMCM_LOCKED_OFFSET 0
`define WB_FMC_250M_4CH_CSR_FMC_STA_MMCM_LOCKED 32'h00000001
`define WB_FMC_250M_4CH_CSR_FMC_STA_PWR_GOOD_OFFSET 1
`define WB_FMC_250M_4CH_CSR_FMC_STA_PWR_GOOD 32'h00000002
`define WB_FMC_250M_4CH_CSR_FMC_STA_PRST_OFFSET 2
`define WB_FMC_250M_4CH_CSR_FMC_STA_PRST 32'h00000004
`define WB_FMC_250M_4CH_CSR_FMC_STA_RESERVED_OFFSET 3
`define WB_FMC_250M_4CH_CSR_FMC_STA_RESERVED 32'h7ffffff8
`define ADDR_WB_FMC_250M_4CH_CSR_CLK_DISTRIB 7'h4
`define WB_FMC_250M_4CH_CSR_CLK_DISTRIB_SI571_OE_OFFSET 0
`define WB_FMC_250M_4CH_CSR_CLK_DISTRIB_SI571_OE 32'h00000001
`define WB_FMC_250M_4CH_CSR_CLK_DISTRIB_PLL_FUNCTION_OFFSET 1
`define WB_FMC_250M_4CH_CSR_CLK_DISTRIB_PLL_FUNCTION 32'h00000002
`define WB_FMC_250M_4CH_CSR_CLK_DISTRIB_PLL_STATUS_OFFSET 2
`define WB_FMC_250M_4CH_CSR_CLK_DISTRIB_PLL_STATUS 32'h00000004
`define WB_FMC_250M_4CH_CSR_CLK_DISTRIB_CLK_SEL_OFFSET 3
`define WB_FMC_250M_4CH_CSR_CLK_DISTRIB_CLK_SEL 32'h00000008
`define WB_FMC_250M_4CH_CSR_CLK_DISTRIB_RESERVED_OFFSET 4
`define WB_FMC_250M_4CH_CSR_CLK_DISTRIB_RESERVED 32'hfffffff0
`define ADDR_WB_FMC_250M_4CH_CSR_MONITOR 7'h8
`define WB_FMC_250M_4CH_CSR_MONITOR_TEST_DATA_EN_OFFSET 0
`define WB_FMC_250M_4CH_CSR_MONITOR_TEST_DATA_EN 32'h00000001
`define WB_FMC_250M_4CH_CSR_MONITOR_LED1_OFFSET 1
`define WB_FMC_250M_4CH_CSR_MONITOR_LED1 32'h00000002
`define WB_FMC_250M_4CH_CSR_MONITOR_LED2_OFFSET 2
`define WB_FMC_250M_4CH_CSR_MONITOR_LED2 32'h00000004
`define WB_FMC_250M_4CH_CSR_MONITOR_LED3_OFFSET 3
`define WB_FMC_250M_4CH_CSR_MONITOR_LED3 32'h00000008
`define WB_FMC_250M_4CH_CSR_MONITOR_MON_DEV_OFFSET 4
`define WB_FMC_250M_4CH_CSR_MONITOR_MON_DEV 32'h00000010
`define WB_FMC_250M_4CH_CSR_MONITOR_RESERVED_OFFSET 5
`define WB_FMC_250M_4CH_CSR_MONITOR_RESERVED 32'hffffffe0
`define ADDR_WB_FMC_250M_4CH_CSR_TRIGGER 7'hc
`define WB_FMC_250M_4CH_CSR_TRIGGER_DIR_OFFSET 0
`define WB_FMC_250M_4CH_CSR_TRIGGER_DIR 32'h00000001
`define WB_FMC_250M_4CH_CSR_TRIGGER_TERM_OFFSET 1
`define WB_FMC_250M_4CH_CSR_TRIGGER_TERM 32'h00000002
`define WB_FMC_250M_4CH_CSR_TRIGGER_TRIG_VAL_OFFSET 2
`define WB_FMC_250M_4CH_CSR_TRIGGER_TRIG_VAL 32'h00000004
`define WB_FMC_250M_4CH_CSR_TRIGGER_RESERVED_OFFSET 3
`define WB_FMC_250M_4CH_CSR_TRIGGER_RESERVED 32'hfffffff8
`define ADDR_WB_FMC_250M_4CH_CSR_ADC_STA 7'h10
`define WB_FMC_250M_4CH_CSR_ADC_STA_CLK_CHAINS_OFFSET 0
`define WB_FMC_250M_4CH_CSR_ADC_STA_CLK_CHAINS 32'h0000000f
`define WB_FMC_250M_4CH_CSR_ADC_STA_RESERVED_CLK_CHAINS_OFFSET 4
`define WB_FMC_250M_4CH_CSR_ADC_STA_RESERVED_CLK_CHAINS 32'h000000f0
`define WB_FMC_250M_4CH_CSR_ADC_STA_DATA_CHAINS_OFFSET 8
`define WB_FMC_250M_4CH_CSR_ADC_STA_DATA_CHAINS 32'h00000f00
`define WB_FMC_250M_4CH_CSR_ADC_STA_RESERVED_DATA_CHAINS_OFFSET 12
`define WB_FMC_250M_4CH_CSR_ADC_STA_RESERVED_DATA_CHAINS 32'h0000f000
`define WB_FMC_250M_4CH_CSR_ADC_STA_ADC_PKT_SIZE_OFFSET 16
`define WB_FMC_250M_4CH_CSR_ADC_STA_ADC_PKT_SIZE 32'hffff0000
`define ADDR_WB_FMC_250M_4CH_CSR_ADC_CTL 7'h14
`define WB_FMC_250M_4CH_CSR_ADC_CTL_UPDATE_CLK_DLY_OFFSET 0
`define WB_FMC_250M_4CH_CSR_ADC_CTL_UPDATE_CLK_DLY 32'h00000001
`define WB_FMC_250M_4CH_CSR_ADC_CTL_UPDATE_DATA_DLY_OFFSET 1
`define WB_FMC_250M_4CH_CSR_ADC_CTL_UPDATE_DATA_DLY 32'h00000002
`define WB_FMC_250M_4CH_CSR_ADC_CTL_RST_ADCS_OFFSET 2
`define WB_FMC_250M_4CH_CSR_ADC_CTL_RST_ADCS 32'h00000004
`define WB_FMC_250M_4CH_CSR_ADC_CTL_RST_DIV_ADCS_OFFSET 3
`define WB_FMC_250M_4CH_CSR_ADC_CTL_RST_DIV_ADCS 32'h00000008
`define WB_FMC_250M_4CH_CSR_ADC_CTL_RESERVED_OFFSET 4
`define WB_FMC_250M_4CH_CSR_ADC_CTL_RESERVED 32'hfffffff0
`define ADDR_WB_FMC_250M_4CH_CSR_CH0_STA 7'h18
`define WB_FMC_250M_4CH_CSR_CH0_STA_VAL_OFFSET 0
`define WB_FMC_250M_4CH_CSR_CH0_STA_VAL 32'h0000ffff
`define WB_FMC_250M_4CH_CSR_CH0_STA_RESERVED_OFFSET 16
`define WB_FMC_250M_4CH_CSR_CH0_STA_RESERVED 32'hffff0000
`define ADDR_WB_FMC_250M_4CH_CSR_CH0_FN_DLY 7'h1c
`define WB_FMC_250M_4CH_CSR_CH0_FN_DLY_CLK_CHAIN_DLY_OFFSET 0
`define WB_FMC_250M_4CH_CSR_CH0_FN_DLY_CLK_CHAIN_DLY 32'h0000001f
`define WB_FMC_250M_4CH_CSR_CH0_FN_DLY_RESERVED_CLK_CHAIN_DLY_OFFSET 5
`define WB_FMC_250M_4CH_CSR_CH0_FN_DLY_RESERVED_CLK_CHAIN_DLY 32'h000000e0
`define WB_FMC_250M_4CH_CSR_CH0_FN_DLY_DATA_CHAIN_DLY_OFFSET 8
`define WB_FMC_250M_4CH_CSR_CH0_FN_DLY_DATA_CHAIN_DLY 32'h00001f00
`define WB_FMC_250M_4CH_CSR_CH0_FN_DLY_RESERVED_DATA_CHAIN_DLY_OFFSET 13
`define WB_FMC_250M_4CH_CSR_CH0_FN_DLY_RESERVED_DATA_CHAIN_DLY 32'h0000e000
`define WB_FMC_250M_4CH_CSR_CH0_FN_DLY_INC_CLK_CHAIN_DLY_OFFSET 16
`define WB_FMC_250M_4CH_CSR_CH0_FN_DLY_INC_CLK_CHAIN_DLY 32'h00010000
`define WB_FMC_250M_4CH_CSR_CH0_FN_DLY_DEC_CLK_CHAIN_DLY_OFFSET 17
`define WB_FMC_250M_4CH_CSR_CH0_FN_DLY_DEC_CLK_CHAIN_DLY 32'h00020000
`define WB_FMC_250M_4CH_CSR_CH0_FN_DLY_RESERVED_CLK_INCDEC_DLY_OFFSET 18
`define WB_FMC_250M_4CH_CSR_CH0_FN_DLY_RESERVED_CLK_INCDEC_DLY 32'h00fc0000
`define WB_FMC_250M_4CH_CSR_CH0_FN_DLY_INC_DATA_CHAIN_DLY_OFFSET 24
`define WB_FMC_250M_4CH_CSR_CH0_FN_DLY_INC_DATA_CHAIN_DLY 32'h01000000
`define WB_FMC_250M_4CH_CSR_CH0_FN_DLY_DEC_DATA_CHAIN_DLY_OFFSET 25
`define WB_FMC_250M_4CH_CSR_CH0_FN_DLY_DEC_DATA_CHAIN_DLY 32'h02000000
`define WB_FMC_250M_4CH_CSR_CH0_FN_DLY_RESERVED_DATA_INCDEC_DLY_OFFSET 26
`define WB_FMC_250M_4CH_CSR_CH0_FN_DLY_RESERVED_DATA_INCDEC_DLY 32'hfc000000
`define ADDR_WB_FMC_250M_4CH_CSR_CH0_CS_DLY 7'h20
`define WB_FMC_250M_4CH_CSR_CH0_CS_DLY_FE_DLY_OFFSET 0
`define WB_FMC_250M_4CH_CSR_CH0_CS_DLY_FE_DLY 32'h00000003
`define WB_FMC_250M_4CH_CSR_CH0_CS_DLY_RESERVED_FE_DLY_OFFSET 2
`define WB_FMC_250M_4CH_CSR_CH0_CS_DLY_RESERVED_FE_DLY 32'h000000fc
`define WB_FMC_250M_4CH_CSR_CH0_CS_DLY_RG_DLY_OFFSET 8
`define WB_FMC_250M_4CH_CSR_CH0_CS_DLY_RG_DLY 32'h00000300
`define WB_FMC_250M_4CH_CSR_CH0_CS_DLY_RESERVED_RG_DLY_OFFSET 10
`define WB_FMC_250M_4CH_CSR_CH0_CS_DLY_RESERVED_RG_DLY 32'hfffffc00
`define ADDR_WB_FMC_250M_4CH_CSR_CH1_STA 7'h24
`define WB_FMC_250M_4CH_CSR_CH1_STA_VAL_OFFSET 0
`define WB_FMC_250M_4CH_CSR_CH1_STA_VAL 32'h0000ffff
`define WB_FMC_250M_4CH_CSR_CH1_STA_RESERVED_OFFSET 16
`define WB_FMC_250M_4CH_CSR_CH1_STA_RESERVED 32'hffff0000
`define ADDR_WB_FMC_250M_4CH_CSR_CH1_FN_DLY 7'h28
`define WB_FMC_250M_4CH_CSR_CH1_FN_DLY_CLK_CHAIN_DLY_OFFSET 0
`define WB_FMC_250M_4CH_CSR_CH1_FN_DLY_CLK_CHAIN_DLY 32'h0000001f
`define WB_FMC_250M_4CH_CSR_CH1_FN_DLY_RESERVED_CLK_CHAIN_DLY_OFFSET 5
`define WB_FMC_250M_4CH_CSR_CH1_FN_DLY_RESERVED_CLK_CHAIN_DLY 32'h000000e0
`define WB_FMC_250M_4CH_CSR_CH1_FN_DLY_DATA_CHAIN_DLY_OFFSET 8
`define WB_FMC_250M_4CH_CSR_CH1_FN_DLY_DATA_CHAIN_DLY 32'h00001f00
`define WB_FMC_250M_4CH_CSR_CH1_FN_DLY_RESERVED_DATA_CHAIN_DLY_OFFSET 13
`define WB_FMC_250M_4CH_CSR_CH1_FN_DLY_RESERVED_DATA_CHAIN_DLY 32'h0000e000
`define WB_FMC_250M_4CH_CSR_CH1_FN_DLY_INC_CLK_CHAIN_DLY_OFFSET 16
`define WB_FMC_250M_4CH_CSR_CH1_FN_DLY_INC_CLK_CHAIN_DLY 32'h00010000
`define WB_FMC_250M_4CH_CSR_CH1_FN_DLY_DEC_CLK_CHAIN_DLY_OFFSET 17
`define WB_FMC_250M_4CH_CSR_CH1_FN_DLY_DEC_CLK_CHAIN_DLY 32'h00020000
`define WB_FMC_250M_4CH_CSR_CH1_FN_DLY_RESERVED_CLK_INCDEC_DLY_OFFSET 18
`define WB_FMC_250M_4CH_CSR_CH1_FN_DLY_RESERVED_CLK_INCDEC_DLY 32'h00fc0000
`define WB_FMC_250M_4CH_CSR_CH1_FN_DLY_INC_DATA_CHAIN_DLY_OFFSET 24
`define WB_FMC_250M_4CH_CSR_CH1_FN_DLY_INC_DATA_CHAIN_DLY 32'h01000000
`define WB_FMC_250M_4CH_CSR_CH1_FN_DLY_DEC_DATA_CHAIN_DLY_OFFSET 25
`define WB_FMC_250M_4CH_CSR_CH1_FN_DLY_DEC_DATA_CHAIN_DLY 32'h02000000
`define WB_FMC_250M_4CH_CSR_CH1_FN_DLY_RESERVED_DATA_INCDEC_DLY_OFFSET 26
`define WB_FMC_250M_4CH_CSR_CH1_FN_DLY_RESERVED_DATA_INCDEC_DLY 32'hfc000000
`define ADDR_WB_FMC_250M_4CH_CSR_CH1_CS_DLY 7'h2c
`define WB_FMC_250M_4CH_CSR_CH1_CS_DLY_FE_DLY_OFFSET 0
`define WB_FMC_250M_4CH_CSR_CH1_CS_DLY_FE_DLY 32'h00000003
`define WB_FMC_250M_4CH_CSR_CH1_CS_DLY_RESERVED_FE_DLY_OFFSET 2
`define WB_FMC_250M_4CH_CSR_CH1_CS_DLY_RESERVED_FE_DLY 32'h000000fc
`define WB_FMC_250M_4CH_CSR_CH1_CS_DLY_RG_DLY_OFFSET 8
`define WB_FMC_250M_4CH_CSR_CH1_CS_DLY_RG_DLY 32'h00000300
`define WB_FMC_250M_4CH_CSR_CH1_CS_DLY_RESERVED_RG_DLY_OFFSET 10
`define WB_FMC_250M_4CH_CSR_CH1_CS_DLY_RESERVED_RG_DLY 32'hfffffc00
`define ADDR_WB_FMC_250M_4CH_CSR_CH2_STA 7'h30
`define WB_FMC_250M_4CH_CSR_CH2_STA_VAL_OFFSET 0
`define WB_FMC_250M_4CH_CSR_CH2_STA_VAL 32'h0000ffff
`define WB_FMC_250M_4CH_CSR_CH2_STA_RESERVED_OFFSET 16
`define WB_FMC_250M_4CH_CSR_CH2_STA_RESERVED 32'hffff0000
`define ADDR_WB_FMC_250M_4CH_CSR_CH2_FN_DLY 7'h34
`define WB_FMC_250M_4CH_CSR_CH2_FN_DLY_CLK_CHAIN_DLY_OFFSET 0
`define WB_FMC_250M_4CH_CSR_CH2_FN_DLY_CLK_CHAIN_DLY 32'h0000001f
`define WB_FMC_250M_4CH_CSR_CH2_FN_DLY_RESERVED_CLK_CHAIN_DLY_OFFSET 5
`define WB_FMC_250M_4CH_CSR_CH2_FN_DLY_RESERVED_CLK_CHAIN_DLY 32'h000000e0
`define WB_FMC_250M_4CH_CSR_CH2_FN_DLY_DATA_CHAIN_DLY_OFFSET 8
`define WB_FMC_250M_4CH_CSR_CH2_FN_DLY_DATA_CHAIN_DLY 32'h00001f00
`define WB_FMC_250M_4CH_CSR_CH2_FN_DLY_RESERVED_DATA_CHAIN_DLY_OFFSET 13
`define WB_FMC_250M_4CH_CSR_CH2_FN_DLY_RESERVED_DATA_CHAIN_DLY 32'h0000e000
`define WB_FMC_250M_4CH_CSR_CH2_FN_DLY_INC_CLK_CHAIN_DLY_OFFSET 16
`define WB_FMC_250M_4CH_CSR_CH2_FN_DLY_INC_CLK_CHAIN_DLY 32'h00010000
`define WB_FMC_250M_4CH_CSR_CH2_FN_DLY_DEC_CLK_CHAIN_DLY_OFFSET 17
`define WB_FMC_250M_4CH_CSR_CH2_FN_DLY_DEC_CLK_CHAIN_DLY 32'h00020000
`define WB_FMC_250M_4CH_CSR_CH2_FN_DLY_RESERVED_CLK_INCDEC_DLY_OFFSET 18
`define WB_FMC_250M_4CH_CSR_CH2_FN_DLY_RESERVED_CLK_INCDEC_DLY 32'h00fc0000
`define WB_FMC_250M_4CH_CSR_CH2_FN_DLY_INC_DATA_CHAIN_DLY_OFFSET 24
`define WB_FMC_250M_4CH_CSR_CH2_FN_DLY_INC_DATA_CHAIN_DLY 32'h01000000
`define WB_FMC_250M_4CH_CSR_CH2_FN_DLY_DEC_DATA_CHAIN_DLY_OFFSET 25
`define WB_FMC_250M_4CH_CSR_CH2_FN_DLY_DEC_DATA_CHAIN_DLY 32'h02000000
`define WB_FMC_250M_4CH_CSR_CH2_FN_DLY_RESERVED_DATA_INCDEC_DLY_OFFSET 26
`define WB_FMC_250M_4CH_CSR_CH2_FN_DLY_RESERVED_DATA_INCDEC_DLY 32'hfc000000
`define ADDR_WB_FMC_250M_4CH_CSR_CH2_CS_DLY 7'h38
`define WB_FMC_250M_4CH_CSR_CH2_CS_DLY_FE_DLY_OFFSET 0
`define WB_FMC_250M_4CH_CSR_CH2_CS_DLY_FE_DLY 32'h00000003
`define WB_FMC_250M_4CH_CSR_CH2_CS_DLY_RESERVED_FE_DLY_OFFSET 2
`define WB_FMC_250M_4CH_CSR_CH2_CS_DLY_RESERVED_FE_DLY 32'h000000fc
`define WB_FMC_250M_4CH_CSR_CH2_CS_DLY_RG_DLY_OFFSET 8
`define WB_FMC_250M_4CH_CSR_CH2_CS_DLY_RG_DLY 32'h00000300
`define WB_FMC_250M_4CH_CSR_CH2_CS_DLY_RESERVED_RG_DLY_OFFSET 10
`define WB_FMC_250M_4CH_CSR_CH2_CS_DLY_RESERVED_RG_DLY 32'hfffffc00
`define ADDR_WB_FMC_250M_4CH_CSR_CH3_STA 7'h3c
`define WB_FMC_250M_4CH_CSR_CH3_STA_VAL_OFFSET 0
`define WB_FMC_250M_4CH_CSR_CH3_STA_VAL 32'h0000ffff
`define WB_FMC_250M_4CH_CSR_CH3_STA_RESERVED_OFFSET 16
`define WB_FMC_250M_4CH_CSR_CH3_STA_RESERVED 32'hffff0000
`define ADDR_WB_FMC_250M_4CH_CSR_CH3_FN_DLY 7'h40
`define WB_FMC_250M_4CH_CSR_CH3_FN_DLY_CLK_CHAIN_DLY_OFFSET 0
`define WB_FMC_250M_4CH_CSR_CH3_FN_DLY_CLK_CHAIN_DLY 32'h0000001f
`define WB_FMC_250M_4CH_CSR_CH3_FN_DLY_RESERVED_CLK_CHAIN_DLY_OFFSET 5
`define WB_FMC_250M_4CH_CSR_CH3_FN_DLY_RESERVED_CLK_CHAIN_DLY 32'h000000e0
`define WB_FMC_250M_4CH_CSR_CH3_FN_DLY_DATA_CHAIN_DLY_OFFSET 8
`define WB_FMC_250M_4CH_CSR_CH3_FN_DLY_DATA_CHAIN_DLY 32'h00001f00
`define WB_FMC_250M_4CH_CSR_CH3_FN_DLY_RESERVED_DATA_CHAIN_DLY_OFFSET 13
`define WB_FMC_250M_4CH_CSR_CH3_FN_DLY_RESERVED_DATA_CHAIN_DLY 32'h0000e000
`define WB_FMC_250M_4CH_CSR_CH3_FN_DLY_INC_CLK_CHAIN_DLY_OFFSET 16
`define WB_FMC_250M_4CH_CSR_CH3_FN_DLY_INC_CLK_CHAIN_DLY 32'h00010000
`define WB_FMC_250M_4CH_CSR_CH3_FN_DLY_DEC_CLK_CHAIN_DLY_OFFSET 17
`define WB_FMC_250M_4CH_CSR_CH3_FN_DLY_DEC_CLK_CHAIN_DLY 32'h00020000
`define WB_FMC_250M_4CH_CSR_CH3_FN_DLY_RESERVED_CLK_INCDEC_DLY_OFFSET 18
`define WB_FMC_250M_4CH_CSR_CH3_FN_DLY_RESERVED_CLK_INCDEC_DLY 32'h00fc0000
`define WB_FMC_250M_4CH_CSR_CH3_FN_DLY_INC_DATA_CHAIN_DLY_OFFSET 24
`define WB_FMC_250M_4CH_CSR_CH3_FN_DLY_INC_DATA_CHAIN_DLY 32'h01000000
`define WB_FMC_250M_4CH_CSR_CH3_FN_DLY_DEC_DATA_CHAIN_DLY_OFFSET 25
`define WB_FMC_250M_4CH_CSR_CH3_FN_DLY_DEC_DATA_CHAIN_DLY 32'h02000000
`define WB_FMC_250M_4CH_CSR_CH3_FN_DLY_RESERVED_DATA_INCDEC_DLY_OFFSET 26
`define WB_FMC_250M_4CH_CSR_CH3_FN_DLY_RESERVED_DATA_INCDEC_DLY 32'hfc000000
`define ADDR_WB_FMC_250M_4CH_CSR_CH3_CS_DLY 7'h44
`define WB_FMC_250M_4CH_CSR_CH3_CS_DLY_FE_DLY_OFFSET 0
`define WB_FMC_250M_4CH_CSR_CH3_CS_DLY_FE_DLY 32'h00000003
`define WB_FMC_250M_4CH_CSR_CH3_CS_DLY_RESERVED_FE_DLY_OFFSET 2
`define WB_FMC_250M_4CH_CSR_CH3_CS_DLY_RESERVED_FE_DLY 32'h000000fc
`define WB_FMC_250M_4CH_CSR_CH3_CS_DLY_RG_DLY_OFFSET 8
`define WB_FMC_250M_4CH_CSR_CH3_CS_DLY_RG_DLY 32'h00000300
`define WB_FMC_250M_4CH_CSR_CH3_CS_DLY_RESERVED_RG_DLY_OFFSET 10
`define WB_FMC_250M_4CH_CSR_CH3_CS_DLY_RESERVED_RG_DLY 32'hfffffc00
