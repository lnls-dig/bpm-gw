`define ADDR_DATA_SRC_B2C_R0           3'h0
`define DATA_SRC_B2C_R0_DATA_OFFSET 0
`define DATA_SRC_B2C_R0_DATA 32'hffffffff
`define ADDR_DATA_SRC_B2C_CSR          3'h4
`define DATA_SRC_B2C_CSR_FULL_OFFSET 16
`define DATA_SRC_B2C_CSR_FULL 32'h00010000
`define DATA_SRC_B2C_CSR_EMPTY_OFFSET 17
`define DATA_SRC_B2C_CSR_EMPTY 32'h00020000
`define DATA_SRC_B2C_CSR_USEDW_OFFSET 0
`define DATA_SRC_B2C_CSR_USEDW 32'h000000ff
