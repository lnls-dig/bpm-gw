`define ADDR_WB_FMC_ACTIVE_CLK_CSR_CLK_DISTRIB 2'h0
`define WB_FMC_ACTIVE_CLK_CSR_CLK_DISTRIB_SI571_OE_OFFSET 0
`define WB_FMC_ACTIVE_CLK_CSR_CLK_DISTRIB_SI571_OE 32'h00000001
`define WB_FMC_ACTIVE_CLK_CSR_CLK_DISTRIB_PLL_FUNCTION_OFFSET 1
`define WB_FMC_ACTIVE_CLK_CSR_CLK_DISTRIB_PLL_FUNCTION 32'h00000002
`define WB_FMC_ACTIVE_CLK_CSR_CLK_DISTRIB_PLL_STATUS_OFFSET 2
`define WB_FMC_ACTIVE_CLK_CSR_CLK_DISTRIB_PLL_STATUS 32'h00000004
`define WB_FMC_ACTIVE_CLK_CSR_CLK_DISTRIB_CLK_SEL_OFFSET 3
`define WB_FMC_ACTIVE_CLK_CSR_CLK_DISTRIB_CLK_SEL 32'h00000008
`define WB_FMC_ACTIVE_CLK_CSR_CLK_DISTRIB_RESERVED_OFFSET 4
`define WB_FMC_ACTIVE_CLK_CSR_CLK_DISTRIB_RESERVED 32'hfffffff0
