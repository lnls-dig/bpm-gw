`define ADDR_CTL_IFACE_CTL             3'h0
`define CTL_IFACE_CTL_START_OFFSET 0
`define CTL_IFACE_CTL_START 32'h00000001
`define CTL_IFACE_CTL_DONE_OFFSET 1
`define CTL_IFACE_CTL_DONE 32'h00000002
`define CTL_IFACE_CTL_OVF_OFFSET 2
`define CTL_IFACE_CTL_OVF 32'h00000004
`define ADDR_CTL_IFACE_TR_CNTR         3'h4
