package pos_calc_Consts is
  constant POS_CALC_SIZE : Natural := 276;
  constant ADDR_POS_CALC_DS_TBT_THRES : Natural := 16#0#;
  constant POS_CALC_DS_TBT_THRES_VAL_OFFSET : Natural := 0;
  constant POS_CALC_DS_TBT_THRES_RESERVED_OFFSET : Natural := 26;
  constant ADDR_POS_CALC_DS_FOFB_THRES : Natural := 16#4#;
  constant POS_CALC_DS_FOFB_THRES_VAL_OFFSET : Natural := 0;
  constant POS_CALC_DS_FOFB_THRES_RESERVED_OFFSET : Natural := 26;
  constant ADDR_POS_CALC_DS_MONIT_THRES : Natural := 16#8#;
  constant POS_CALC_DS_MONIT_THRES_VAL_OFFSET : Natural := 0;
  constant POS_CALC_DS_MONIT_THRES_RESERVED_OFFSET : Natural := 26;
  constant ADDR_POS_CALC_KX : Natural := 16#c#;
  constant POS_CALC_KX_VAL_OFFSET : Natural := 0;
  constant POS_CALC_KX_RESERVED_OFFSET : Natural := 25;
  constant ADDR_POS_CALC_KY : Natural := 16#10#;
  constant POS_CALC_KY_VAL_OFFSET : Natural := 0;
  constant POS_CALC_KY_RESERVED_OFFSET : Natural := 25;
  constant ADDR_POS_CALC_KSUM : Natural := 16#14#;
  constant POS_CALC_KSUM_VAL_OFFSET : Natural := 0;
  constant POS_CALC_KSUM_RESERVED_OFFSET : Natural := 25;
  constant ADDR_POS_CALC_DSP_CTNR_TBT : Natural := 16#18#;
  constant POS_CALC_DSP_CTNR_TBT_CH01_OFFSET : Natural := 0;
  constant POS_CALC_DSP_CTNR_TBT_CH23_OFFSET : Natural := 16;
  constant ADDR_POS_CALC_DSP_CTNR_FOFB : Natural := 16#1c#;
  constant POS_CALC_DSP_CTNR_FOFB_CH01_OFFSET : Natural := 0;
  constant POS_CALC_DSP_CTNR_FOFB_CH23_OFFSET : Natural := 16;
  constant ADDR_POS_CALC_DSP_CTNR1_MONIT : Natural := 16#20#;
  constant POS_CALC_DSP_CTNR1_MONIT_CIC_OFFSET : Natural := 0;
  constant POS_CALC_DSP_CTNR1_MONIT_CFIR_OFFSET : Natural := 16;
  constant ADDR_POS_CALC_DSP_CTNR2_MONIT : Natural := 16#24#;
  constant POS_CALC_DSP_CTNR2_MONIT_PFIR_OFFSET : Natural := 0;
  constant POS_CALC_DSP_CTNR2_MONIT_FIR_01_OFFSET : Natural := 16;
  constant ADDR_POS_CALC_DSP_ERR_CLR : Natural := 16#28#;
  constant POS_CALC_DSP_ERR_CLR_TBT_OFFSET : Natural := 0;
  constant POS_CALC_DSP_ERR_CLR_FOFB_OFFSET : Natural := 1;
  constant POS_CALC_DSP_ERR_CLR_MONIT_PART1_OFFSET : Natural := 2;
  constant POS_CALC_DSP_ERR_CLR_MONIT_PART2_OFFSET : Natural := 3;
  constant ADDR_POS_CALC_DDS_CFG : Natural := 16#2c#;
  constant POS_CALC_DDS_CFG_VALID_CH0_OFFSET : Natural := 0;
  constant POS_CALC_DDS_CFG_TEST_DATA_OFFSET : Natural := 1;
  constant POS_CALC_DDS_CFG_RESERVED_CH0_OFFSET : Natural := 2;
  constant POS_CALC_DDS_CFG_VALID_CH1_OFFSET : Natural := 8;
  constant POS_CALC_DDS_CFG_RESERVED_CH1_OFFSET : Natural := 9;
  constant POS_CALC_DDS_CFG_VALID_CH2_OFFSET : Natural := 16;
  constant POS_CALC_DDS_CFG_RESERVED_CH2_OFFSET : Natural := 17;
  constant POS_CALC_DDS_CFG_VALID_CH3_OFFSET : Natural := 24;
  constant POS_CALC_DDS_CFG_RESERVED_CH3_OFFSET : Natural := 25;
  constant ADDR_POS_CALC_DDS_PINC_CH0 : Natural := 16#30#;
  constant POS_CALC_DDS_PINC_CH0_VAL_OFFSET : Natural := 0;
  constant POS_CALC_DDS_PINC_CH0_RESERVED_OFFSET : Natural := 30;
  constant ADDR_POS_CALC_DDS_PINC_CH1 : Natural := 16#34#;
  constant POS_CALC_DDS_PINC_CH1_VAL_OFFSET : Natural := 0;
  constant POS_CALC_DDS_PINC_CH1_RESERVED_OFFSET : Natural := 30;
  constant ADDR_POS_CALC_DDS_PINC_CH2 : Natural := 16#38#;
  constant POS_CALC_DDS_PINC_CH2_VAL_OFFSET : Natural := 0;
  constant POS_CALC_DDS_PINC_CH2_RESERVED_OFFSET : Natural := 30;
  constant ADDR_POS_CALC_DDS_PINC_CH3 : Natural := 16#3c#;
  constant POS_CALC_DDS_PINC_CH3_VAL_OFFSET : Natural := 0;
  constant POS_CALC_DDS_PINC_CH3_RESERVED_OFFSET : Natural := 30;
  constant ADDR_POS_CALC_DDS_POFF_CH0 : Natural := 16#40#;
  constant POS_CALC_DDS_POFF_CH0_VAL_OFFSET : Natural := 0;
  constant POS_CALC_DDS_POFF_CH0_RESERVED_OFFSET : Natural := 30;
  constant ADDR_POS_CALC_DDS_POFF_CH1 : Natural := 16#44#;
  constant POS_CALC_DDS_POFF_CH1_VAL_OFFSET : Natural := 0;
  constant POS_CALC_DDS_POFF_CH1_RESERVED_OFFSET : Natural := 30;
  constant ADDR_POS_CALC_DDS_POFF_CH2 : Natural := 16#48#;
  constant POS_CALC_DDS_POFF_CH2_VAL_OFFSET : Natural := 0;
  constant POS_CALC_DDS_POFF_CH2_RESERVED_OFFSET : Natural := 30;
  constant ADDR_POS_CALC_DDS_POFF_CH3 : Natural := 16#4c#;
  constant POS_CALC_DDS_POFF_CH3_VAL_OFFSET : Natural := 0;
  constant POS_CALC_DDS_POFF_CH3_RESERVED_OFFSET : Natural := 30;
  constant ADDR_POS_CALC_DSP_MONIT_AMP_CH0 : Natural := 16#50#;
  constant ADDR_POS_CALC_DSP_MONIT_AMP_CH1 : Natural := 16#54#;
  constant ADDR_POS_CALC_DSP_MONIT_AMP_CH2 : Natural := 16#58#;
  constant ADDR_POS_CALC_DSP_MONIT_AMP_CH3 : Natural := 16#5c#;
  constant ADDR_POS_CALC_DSP_MONIT_POS_X : Natural := 16#60#;
  constant ADDR_POS_CALC_DSP_MONIT_POS_Y : Natural := 16#64#;
  constant ADDR_POS_CALC_DSP_MONIT_POS_Q : Natural := 16#68#;
  constant ADDR_POS_CALC_DSP_MONIT_POS_SUM : Natural := 16#6c#;
  constant ADDR_POS_CALC_DSP_MONIT_UPDT : Natural := 16#70#;
  constant ADDR_POS_CALC_DSP_MONIT1_AMP_CH0 : Natural := 16#74#;
  constant ADDR_POS_CALC_DSP_MONIT1_AMP_CH1 : Natural := 16#78#;
  constant ADDR_POS_CALC_DSP_MONIT1_AMP_CH2 : Natural := 16#7c#;
  constant ADDR_POS_CALC_DSP_MONIT1_AMP_CH3 : Natural := 16#80#;
  constant ADDR_POS_CALC_DSP_MONIT1_POS_X : Natural := 16#84#;
  constant ADDR_POS_CALC_DSP_MONIT1_POS_Y : Natural := 16#88#;
  constant ADDR_POS_CALC_DSP_MONIT1_POS_Q : Natural := 16#8c#;
  constant ADDR_POS_CALC_DSP_MONIT1_POS_SUM : Natural := 16#90#;
  constant ADDR_POS_CALC_DSP_MONIT1_UPDT : Natural := 16#94#;
  constant ADDR_POS_CALC_AMPFIFO_MONIT : Natural := 16#98#;
  constant POS_CALC_AMPFIFO_MONIT_SIZE : Natural := 20;
  constant ADDR_POS_CALC_AMPFIFO_MONIT_AMPFIFO_MONIT_R0 : Natural := 16#98#;
  constant POS_CALC_AMPFIFO_MONIT_AMPFIFO_MONIT_R0_AMP_CH0_OFFSET : Natural := 0;
  constant ADDR_POS_CALC_AMPFIFO_MONIT_AMPFIFO_MONIT_R1 : Natural := 16#9c#;
  constant POS_CALC_AMPFIFO_MONIT_AMPFIFO_MONIT_R1_AMP_CH1_OFFSET : Natural := 0;
  constant ADDR_POS_CALC_AMPFIFO_MONIT_AMPFIFO_MONIT_R2 : Natural := 16#a0#;
  constant POS_CALC_AMPFIFO_MONIT_AMPFIFO_MONIT_R2_AMP_CH2_OFFSET : Natural := 0;
  constant ADDR_POS_CALC_AMPFIFO_MONIT_AMPFIFO_MONIT_R3 : Natural := 16#a4#;
  constant POS_CALC_AMPFIFO_MONIT_AMPFIFO_MONIT_R3_AMP_CH3_OFFSET : Natural := 0;
  constant ADDR_POS_CALC_AMPFIFO_MONIT_AMPFIFO_MONIT_CSR : Natural := 16#a8#;
  constant POS_CALC_AMPFIFO_MONIT_AMPFIFO_MONIT_CSR_FULL_OFFSET : Natural := 16;
  constant POS_CALC_AMPFIFO_MONIT_AMPFIFO_MONIT_CSR_EMPTY_OFFSET : Natural := 17;
  constant POS_CALC_AMPFIFO_MONIT_AMPFIFO_MONIT_CSR_COUNT_OFFSET : Natural := 0;
  constant ADDR_POS_CALC_POSFIFO_MONIT : Natural := 16#ac#;
  constant POS_CALC_POSFIFO_MONIT_SIZE : Natural := 20;
  constant ADDR_POS_CALC_POSFIFO_MONIT_POSFIFO_MONIT_R0 : Natural := 16#ac#;
  constant POS_CALC_POSFIFO_MONIT_POSFIFO_MONIT_R0_POS_X_OFFSET : Natural := 0;
  constant ADDR_POS_CALC_POSFIFO_MONIT_POSFIFO_MONIT_R1 : Natural := 16#b0#;
  constant POS_CALC_POSFIFO_MONIT_POSFIFO_MONIT_R1_POS_Y_OFFSET : Natural := 0;
  constant ADDR_POS_CALC_POSFIFO_MONIT_POSFIFO_MONIT_R2 : Natural := 16#b4#;
  constant POS_CALC_POSFIFO_MONIT_POSFIFO_MONIT_R2_POS_Q_OFFSET : Natural := 0;
  constant ADDR_POS_CALC_POSFIFO_MONIT_POSFIFO_MONIT_R3 : Natural := 16#b8#;
  constant POS_CALC_POSFIFO_MONIT_POSFIFO_MONIT_R3_POS_SUM_OFFSET : Natural := 0;
  constant ADDR_POS_CALC_POSFIFO_MONIT_POSFIFO_MONIT_CSR : Natural := 16#bc#;
  constant POS_CALC_POSFIFO_MONIT_POSFIFO_MONIT_CSR_FULL_OFFSET : Natural := 16;
  constant POS_CALC_POSFIFO_MONIT_POSFIFO_MONIT_CSR_EMPTY_OFFSET : Natural := 17;
  constant POS_CALC_POSFIFO_MONIT_POSFIFO_MONIT_CSR_COUNT_OFFSET : Natural := 0;
  constant ADDR_POS_CALC_AMPFIFO_MONIT1 : Natural := 16#c0#;
  constant POS_CALC_AMPFIFO_MONIT1_SIZE : Natural := 20;
  constant ADDR_POS_CALC_AMPFIFO_MONIT1_AMPFIFO_MONIT1_R0 : Natural := 16#c0#;
  constant POS_CALC_AMPFIFO_MONIT1_AMPFIFO_MONIT1_R0_AMP_CH0_OFFSET : Natural := 0;
  constant ADDR_POS_CALC_AMPFIFO_MONIT1_AMPFIFO_MONIT1_R1 : Natural := 16#c4#;
  constant POS_CALC_AMPFIFO_MONIT1_AMPFIFO_MONIT1_R1_AMP_CH1_OFFSET : Natural := 0;
  constant ADDR_POS_CALC_AMPFIFO_MONIT1_AMPFIFO_MONIT1_R2 : Natural := 16#c8#;
  constant POS_CALC_AMPFIFO_MONIT1_AMPFIFO_MONIT1_R2_AMP_CH2_OFFSET : Natural := 0;
  constant ADDR_POS_CALC_AMPFIFO_MONIT1_AMPFIFO_MONIT1_R3 : Natural := 16#cc#;
  constant POS_CALC_AMPFIFO_MONIT1_AMPFIFO_MONIT1_R3_AMP_CH3_OFFSET : Natural := 0;
  constant ADDR_POS_CALC_AMPFIFO_MONIT1_AMPFIFO_MONIT1_CSR : Natural := 16#d0#;
  constant POS_CALC_AMPFIFO_MONIT1_AMPFIFO_MONIT1_CSR_FULL_OFFSET : Natural := 16;
  constant POS_CALC_AMPFIFO_MONIT1_AMPFIFO_MONIT1_CSR_EMPTY_OFFSET : Natural := 17;
  constant POS_CALC_AMPFIFO_MONIT1_AMPFIFO_MONIT1_CSR_COUNT_OFFSET : Natural := 0;
  constant ADDR_POS_CALC_POSFIFO_MONIT1 : Natural := 16#d4#;
  constant POS_CALC_POSFIFO_MONIT1_SIZE : Natural := 20;
  constant ADDR_POS_CALC_POSFIFO_MONIT1_POSFIFO_MONIT1_R0 : Natural := 16#d4#;
  constant POS_CALC_POSFIFO_MONIT1_POSFIFO_MONIT1_R0_POS_X_OFFSET : Natural := 0;
  constant ADDR_POS_CALC_POSFIFO_MONIT1_POSFIFO_MONIT1_R1 : Natural := 16#d8#;
  constant POS_CALC_POSFIFO_MONIT1_POSFIFO_MONIT1_R1_POS_Y_OFFSET : Natural := 0;
  constant ADDR_POS_CALC_POSFIFO_MONIT1_POSFIFO_MONIT1_R2 : Natural := 16#dc#;
  constant POS_CALC_POSFIFO_MONIT1_POSFIFO_MONIT1_R2_POS_Q_OFFSET : Natural := 0;
  constant ADDR_POS_CALC_POSFIFO_MONIT1_POSFIFO_MONIT1_R3 : Natural := 16#e0#;
  constant POS_CALC_POSFIFO_MONIT1_POSFIFO_MONIT1_R3_POS_SUM_OFFSET : Natural := 0;
  constant ADDR_POS_CALC_POSFIFO_MONIT1_POSFIFO_MONIT1_CSR : Natural := 16#e4#;
  constant POS_CALC_POSFIFO_MONIT1_POSFIFO_MONIT1_CSR_FULL_OFFSET : Natural := 16;
  constant POS_CALC_POSFIFO_MONIT1_POSFIFO_MONIT1_CSR_EMPTY_OFFSET : Natural := 17;
  constant POS_CALC_POSFIFO_MONIT1_POSFIFO_MONIT1_CSR_COUNT_OFFSET : Natural := 0;
  constant ADDR_POS_CALC_SW_TAG : Natural := 16#e8#;
  constant POS_CALC_SW_TAG_EN_OFFSET : Natural := 0;
  constant POS_CALC_SW_TAG_DESYNC_CNT_RST_OFFSET : Natural := 8;
  constant POS_CALC_SW_TAG_DESYNC_CNT_OFFSET : Natural := 9;
  constant ADDR_POS_CALC_SW_DATA_MASK : Natural := 16#ec#;
  constant POS_CALC_SW_DATA_MASK_EN_OFFSET : Natural := 0;
  constant POS_CALC_SW_DATA_MASK_SAMPLES_OFFSET : Natural := 1;
  constant ADDR_POS_CALC_TBT_TAG : Natural := 16#f0#;
  constant POS_CALC_TBT_TAG_EN_OFFSET : Natural := 0;
  constant POS_CALC_TBT_TAG_DLY_OFFSET : Natural := 1;
  constant POS_CALC_TBT_TAG_DESYNC_CNT_RST_OFFSET : Natural := 17;
  constant POS_CALC_TBT_TAG_DESYNC_CNT_OFFSET : Natural := 18;
  constant ADDR_POS_CALC_TBT_DATA_MASK_CTL : Natural := 16#f4#;
  constant POS_CALC_TBT_DATA_MASK_CTL_EN_OFFSET : Natural := 0;
  constant ADDR_POS_CALC_TBT_DATA_MASK_SAMPLES : Natural := 16#f8#;
  constant POS_CALC_TBT_DATA_MASK_SAMPLES_BEG_OFFSET : Natural := 0;
  constant POS_CALC_TBT_DATA_MASK_SAMPLES_END_OFFSET : Natural := 16;
  constant ADDR_POS_CALC_MONIT1_TAG : Natural := 16#fc#;
  constant POS_CALC_MONIT1_TAG_EN_OFFSET : Natural := 0;
  constant POS_CALC_MONIT1_TAG_DLY_OFFSET : Natural := 1;
  constant POS_CALC_MONIT1_TAG_DESYNC_CNT_RST_OFFSET : Natural := 17;
  constant POS_CALC_MONIT1_TAG_DESYNC_CNT_OFFSET : Natural := 18;
  constant ADDR_POS_CALC_MONIT1_DATA_MASK_CTL : Natural := 16#100#;
  constant POS_CALC_MONIT1_DATA_MASK_CTL_EN_OFFSET : Natural := 0;
  constant ADDR_POS_CALC_MONIT1_DATA_MASK_SAMPLES : Natural := 16#104#;
  constant POS_CALC_MONIT1_DATA_MASK_SAMPLES_BEG_OFFSET : Natural := 0;
  constant POS_CALC_MONIT1_DATA_MASK_SAMPLES_END_OFFSET : Natural := 16;
  constant ADDR_POS_CALC_MONIT_TAG : Natural := 16#108#;
  constant POS_CALC_MONIT_TAG_EN_OFFSET : Natural := 0;
  constant POS_CALC_MONIT_TAG_DLY_OFFSET : Natural := 1;
  constant POS_CALC_MONIT_TAG_DESYNC_CNT_RST_OFFSET : Natural := 17;
  constant POS_CALC_MONIT_TAG_DESYNC_CNT_OFFSET : Natural := 18;
  constant ADDR_POS_CALC_MONIT_DATA_MASK_CTL : Natural := 16#10c#;
  constant POS_CALC_MONIT_DATA_MASK_CTL_EN_OFFSET : Natural := 0;
  constant ADDR_POS_CALC_MONIT_DATA_MASK_SAMPLES : Natural := 16#110#;
  constant POS_CALC_MONIT_DATA_MASK_SAMPLES_BEG_OFFSET : Natural := 0;
  constant POS_CALC_MONIT_DATA_MASK_SAMPLES_END_OFFSET : Natural := 16;
end package pos_calc_Consts;
