`define ADDR_FMC516_FMC_STA            7'h0
`define FMC516_FMC_STA_LMK_LOCKED_OFFSET 0
`define FMC516_FMC_STA_LMK_LOCKED 32'h00000001
`define FMC516_FMC_STA_MMCM_LOCKED_OFFSET 1
`define FMC516_FMC_STA_MMCM_LOCKED 32'h00000002
`define FMC516_FMC_STA_PWR_GOOD_OFFSET 2
`define FMC516_FMC_STA_PWR_GOOD 32'h00000004
`define FMC516_FMC_STA_PRST_OFFSET 3
`define FMC516_FMC_STA_PRST 32'h00000008
`define FMC516_FMC_STA_RESERVED_OFFSET 4
`define FMC516_FMC_STA_RESERVED 32'hfffffff0
`define ADDR_FMC516_FMC_CTL            7'h4
`define FMC516_FMC_CTL_TEST_DATA_EN_OFFSET 0
`define FMC516_FMC_CTL_TEST_DATA_EN 32'h00000001
`define FMC516_FMC_CTL_LED_0_OFFSET 1
`define FMC516_FMC_CTL_LED_0 32'h00000002
`define FMC516_FMC_CTL_LED_1_OFFSET 2
`define FMC516_FMC_CTL_LED_1 32'h00000004
`define FMC516_FMC_CTL_CLK_SEL_OFFSET 3
`define FMC516_FMC_CTL_CLK_SEL 32'h00000008
`define FMC516_FMC_CTL_VCXO_OUT_EN_OFFSET 4
`define FMC516_FMC_CTL_VCXO_OUT_EN 32'h00000010
`define FMC516_FMC_CTL_RESERVED_OFFSET 5
`define FMC516_FMC_CTL_RESERVED 32'hffffffe0
`define ADDR_FMC516_TRIG_CFG           7'h8
`define FMC516_TRIG_CFG_HW_TRIG_POL_OFFSET 0
`define FMC516_TRIG_CFG_HW_TRIG_POL 32'h00000001
`define FMC516_TRIG_CFG_HW_TRIG_EN_OFFSET 1
`define FMC516_TRIG_CFG_HW_TRIG_EN 32'h00000002
`define FMC516_TRIG_CFG_RESERVED_OFFSET 2
`define FMC516_TRIG_CFG_RESERVED 32'hfffffffc
`define ADDR_FMC516_ADC_STA            7'hc
`define FMC516_ADC_STA_CLK_CHAINS_OFFSET 0
`define FMC516_ADC_STA_CLK_CHAINS 32'h0000000f
`define FMC516_ADC_STA_RESERVED_CLK_CHAINS_OFFSET 4
`define FMC516_ADC_STA_RESERVED_CLK_CHAINS 32'h000000f0
`define FMC516_ADC_STA_DATA_CHAINS_OFFSET 8
`define FMC516_ADC_STA_DATA_CHAINS 32'h00000f00
`define FMC516_ADC_STA_RESERVED_DATA_CHAINS_OFFSET 12
`define FMC516_ADC_STA_RESERVED_DATA_CHAINS 32'h0000f000
`define FMC516_ADC_STA_ADC_PKT_SIZE_OFFSET 16
`define FMC516_ADC_STA_ADC_PKT_SIZE 32'hffff0000
`define ADDR_FMC516_ADC_CTL            7'h10
`define FMC516_ADC_CTL_UPDATE_CLK_DLY_OFFSET 0
`define FMC516_ADC_CTL_UPDATE_CLK_DLY 32'h00000001
`define FMC516_ADC_CTL_UPDATE_DATA_DLY_OFFSET 1
`define FMC516_ADC_CTL_UPDATE_DATA_DLY 32'h00000002
`define FMC516_ADC_CTL_RST_ADCS_OFFSET 2
`define FMC516_ADC_CTL_RST_ADCS 32'h00000004
`define FMC516_ADC_CTL_RST_DIV_ADCS_OFFSET 3
`define FMC516_ADC_CTL_RST_DIV_ADCS 32'h00000008
`define FMC516_ADC_CTL_RESERVED_OFFSET 4
`define FMC516_ADC_CTL_RESERVED 32'hfffffff0
`define ADDR_FMC516_CH0_STA            7'h14
`define FMC516_CH0_STA_VAL_OFFSET 0
`define FMC516_CH0_STA_VAL 32'h0000ffff
`define FMC516_CH0_STA_RESERVED_OFFSET 16
`define FMC516_CH0_STA_RESERVED 32'hffff0000
`define ADDR_FMC516_CH0_CTL            7'h18
`define FMC516_CH0_CTL_CLK_CHAIN_DLY_OFFSET 0
`define FMC516_CH0_CTL_CLK_CHAIN_DLY 32'h0000001f
`define FMC516_CH0_CTL_RESERVED_CLK_CHAIN_DLY_OFFSET 5
`define FMC516_CH0_CTL_RESERVED_CLK_CHAIN_DLY 32'h000000e0
`define FMC516_CH0_CTL_DATA_CHAIN_DLY_OFFSET 8
`define FMC516_CH0_CTL_DATA_CHAIN_DLY 32'h00001f00
`define FMC516_CH0_CTL_RESERVED_DATA_CHAIN_DLY_OFFSET 13
`define FMC516_CH0_CTL_RESERVED_DATA_CHAIN_DLY 32'h0000e000
`define FMC516_CH0_CTL_INC_CLK_CHAIN_DLY_OFFSET 16
`define FMC516_CH0_CTL_INC_CLK_CHAIN_DLY 32'h00010000
`define FMC516_CH0_CTL_DEC_CLK_CHAIN_DLY_OFFSET 17
`define FMC516_CH0_CTL_DEC_CLK_CHAIN_DLY 32'h00020000
`define FMC516_CH0_CTL_RESERVED_CLK_INCDEC_DLY_OFFSET 18
`define FMC516_CH0_CTL_RESERVED_CLK_INCDEC_DLY 32'h00fc0000
`define FMC516_CH0_CTL_INC_DATA_CHAIN_DLY_OFFSET 24
`define FMC516_CH0_CTL_INC_DATA_CHAIN_DLY 32'h01000000
`define FMC516_CH0_CTL_DEC_DATA_CHAIN_DLY_OFFSET 25
`define FMC516_CH0_CTL_DEC_DATA_CHAIN_DLY 32'h02000000
`define FMC516_CH0_CTL_RESERVED_DATA_INCDEC_DLY_OFFSET 26
`define FMC516_CH0_CTL_RESERVED_DATA_INCDEC_DLY 32'hfc000000
`define ADDR_FMC516_CH0_DLY_CTL        7'h1c
`define FMC516_CH0_DLY_CTL_FE_DLY_OFFSET 0
`define FMC516_CH0_DLY_CTL_FE_DLY 32'h00000003
`define FMC516_CH0_DLY_CTL_RESERVED_FE_DLY_OFFSET 2
`define FMC516_CH0_DLY_CTL_RESERVED_FE_DLY 32'hfffffffc
`define ADDR_FMC516_CH1_STA            7'h20
`define FMC516_CH1_STA_VAL_OFFSET 0
`define FMC516_CH1_STA_VAL 32'h0000ffff
`define FMC516_CH1_STA_RESERVED_OFFSET 16
`define FMC516_CH1_STA_RESERVED 32'hffff0000
`define ADDR_FMC516_CH1_CTL            7'h24
`define FMC516_CH1_CTL_CLK_CHAIN_DLY_OFFSET 0
`define FMC516_CH1_CTL_CLK_CHAIN_DLY 32'h0000001f
`define FMC516_CH1_CTL_RESERVED_CLK_CHAIN_DLY_OFFSET 5
`define FMC516_CH1_CTL_RESERVED_CLK_CHAIN_DLY 32'h000000e0
`define FMC516_CH1_CTL_DATA_CHAIN_DLY_OFFSET 8
`define FMC516_CH1_CTL_DATA_CHAIN_DLY 32'h00001f00
`define FMC516_CH1_CTL_RESERVED_DATA_CHAIN_DLY_OFFSET 13
`define FMC516_CH1_CTL_RESERVED_DATA_CHAIN_DLY 32'h0000e000
`define FMC516_CH1_CTL_INC_CLK_CHAIN_DLY_OFFSET 16
`define FMC516_CH1_CTL_INC_CLK_CHAIN_DLY 32'h00010000
`define FMC516_CH1_CTL_DEC_CLK_CHAIN_DLY_OFFSET 17
`define FMC516_CH1_CTL_DEC_CLK_CHAIN_DLY 32'h00020000
`define FMC516_CH1_CTL_RESERVED_CLK_INCDEC_DLY_OFFSET 18
`define FMC516_CH1_CTL_RESERVED_CLK_INCDEC_DLY 32'h00fc0000
`define FMC516_CH1_CTL_INC_DATA_CHAIN_DLY_OFFSET 24
`define FMC516_CH1_CTL_INC_DATA_CHAIN_DLY 32'h01000000
`define FMC516_CH1_CTL_DEC_DATA_CHAIN_DLY_OFFSET 25
`define FMC516_CH1_CTL_DEC_DATA_CHAIN_DLY 32'h02000000
`define FMC516_CH1_CTL_RESERVED_DATA_INCDEC_DLY_OFFSET 26
`define FMC516_CH1_CTL_RESERVED_DATA_INCDEC_DLY 32'hfc000000
`define ADDR_FMC516_CH1_DLY_CTL        7'h28
`define FMC516_CH1_DLY_CTL_FE_DLY_OFFSET 0
`define FMC516_CH1_DLY_CTL_FE_DLY 32'h00000003
`define FMC516_CH1_DLY_CTL_RESERVED_FE_DLY_OFFSET 2
`define FMC516_CH1_DLY_CTL_RESERVED_FE_DLY 32'hfffffffc
`define ADDR_FMC516_CH2_STA            7'h2c
`define FMC516_CH2_STA_VAL_OFFSET 0
`define FMC516_CH2_STA_VAL 32'h0000ffff
`define FMC516_CH2_STA_RESERVED_OFFSET 16
`define FMC516_CH2_STA_RESERVED 32'hffff0000
`define ADDR_FMC516_CH2_CTL            7'h30
`define FMC516_CH2_CTL_CLK_CHAIN_DLY_OFFSET 0
`define FMC516_CH2_CTL_CLK_CHAIN_DLY 32'h0000001f
`define FMC516_CH2_CTL_RESERVED_CLK_CHAIN_DLY_OFFSET 5
`define FMC516_CH2_CTL_RESERVED_CLK_CHAIN_DLY 32'h000000e0
`define FMC516_CH2_CTL_DATA_CHAIN_DLY_OFFSET 8
`define FMC516_CH2_CTL_DATA_CHAIN_DLY 32'h00001f00
`define FMC516_CH2_CTL_RESERVED_DATA_CHAIN_DLY_OFFSET 13
`define FMC516_CH2_CTL_RESERVED_DATA_CHAIN_DLY 32'h0000e000
`define FMC516_CH2_CTL_INC_CLK_CHAIN_DLY_OFFSET 16
`define FMC516_CH2_CTL_INC_CLK_CHAIN_DLY 32'h00010000
`define FMC516_CH2_CTL_DEC_CLK_CHAIN_DLY_OFFSET 17
`define FMC516_CH2_CTL_DEC_CLK_CHAIN_DLY 32'h00020000
`define FMC516_CH2_CTL_RESERVED_CLK_INCDEC_DLY_OFFSET 18
`define FMC516_CH2_CTL_RESERVED_CLK_INCDEC_DLY 32'h00fc0000
`define FMC516_CH2_CTL_INC_DATA_CHAIN_DLY_OFFSET 24
`define FMC516_CH2_CTL_INC_DATA_CHAIN_DLY 32'h01000000
`define FMC516_CH2_CTL_DEC_DATA_CHAIN_DLY_OFFSET 25
`define FMC516_CH2_CTL_DEC_DATA_CHAIN_DLY 32'h02000000
`define FMC516_CH2_CTL_RESERVED_DATA_INCDEC_DLY_OFFSET 26
`define FMC516_CH2_CTL_RESERVED_DATA_INCDEC_DLY 32'hfc000000
`define ADDR_FMC516_CH2_DLY_CTL        7'h34
`define FMC516_CH2_DLY_CTL_FE_DLY_OFFSET 0
`define FMC516_CH2_DLY_CTL_FE_DLY 32'h00000003
`define FMC516_CH2_DLY_CTL_RESERVED_FE_DLY_OFFSET 2
`define FMC516_CH2_DLY_CTL_RESERVED_FE_DLY 32'hfffffffc
`define ADDR_FMC516_CH3_STA            7'h38
`define FMC516_CH3_STA_VAL_OFFSET 0
`define FMC516_CH3_STA_VAL 32'h0000ffff
`define FMC516_CH3_STA_RESERVED_OFFSET 16
`define FMC516_CH3_STA_RESERVED 32'hffff0000
`define ADDR_FMC516_CH3_CTL            7'h3c
`define FMC516_CH3_CTL_CLK_CHAIN_DLY_OFFSET 0
`define FMC516_CH3_CTL_CLK_CHAIN_DLY 32'h0000001f
`define FMC516_CH3_CTL_RESERVED_CLK_CHAIN_DLY_OFFSET 5
`define FMC516_CH3_CTL_RESERVED_CLK_CHAIN_DLY 32'h000000e0
`define FMC516_CH3_CTL_DATA_CHAIN_DLY_OFFSET 8
`define FMC516_CH3_CTL_DATA_CHAIN_DLY 32'h00001f00
`define FMC516_CH3_CTL_RESERVED_DATA_CHAIN_DLY_OFFSET 13
`define FMC516_CH3_CTL_RESERVED_DATA_CHAIN_DLY 32'h0000e000
`define FMC516_CH3_CTL_INC_CLK_CHAIN_DLY_OFFSET 16
`define FMC516_CH3_CTL_INC_CLK_CHAIN_DLY 32'h00010000
`define FMC516_CH3_CTL_DEC_CLK_CHAIN_DLY_OFFSET 17
`define FMC516_CH3_CTL_DEC_CLK_CHAIN_DLY 32'h00020000
`define FMC516_CH3_CTL_RESERVED_CLK_INCDEC_DLY_OFFSET 18
`define FMC516_CH3_CTL_RESERVED_CLK_INCDEC_DLY 32'h00fc0000
`define FMC516_CH3_CTL_INC_DATA_CHAIN_DLY_OFFSET 24
`define FMC516_CH3_CTL_INC_DATA_CHAIN_DLY 32'h01000000
`define FMC516_CH3_CTL_DEC_DATA_CHAIN_DLY_OFFSET 25
`define FMC516_CH3_CTL_DEC_DATA_CHAIN_DLY 32'h02000000
`define FMC516_CH3_CTL_RESERVED_DATA_INCDEC_DLY_OFFSET 26
`define FMC516_CH3_CTL_RESERVED_DATA_INCDEC_DLY 32'hfc000000
`define ADDR_FMC516_CH3_DLY_CTL        7'h40
`define FMC516_CH3_DLY_CTL_FE_DLY_OFFSET 0
`define FMC516_CH3_DLY_CTL_FE_DLY 32'h00000003
`define FMC516_CH3_DLY_CTL_RESERVED_FE_DLY_OFFSET 2
`define FMC516_CH3_DLY_CTL_RESERVED_FE_DLY 32'hfffffffc
