`define ADDR_DATA_SINK_FIFO_C2B_R0     4'h0
`define DATA_SINK_FIFO_C2B_R0_DATA_OFFSET 0
`define DATA_SINK_FIFO_C2B_R0_DATA 32'hffffffff
`define ADDR_DATA_SINK_FIFO_C2B_R1     4'h4
`define DATA_SINK_FIFO_C2B_R1_LAST_OFFSET 0
`define DATA_SINK_FIFO_C2B_R1_LAST 32'h00000001
`define ADDR_DATA_SINK_FIFO_C2B_CSR    4'h8
`define DATA_SINK_FIFO_C2B_CSR_FULL_OFFSET 16
`define DATA_SINK_FIFO_C2B_CSR_FULL 32'h00010000
`define DATA_SINK_FIFO_C2B_CSR_EMPTY_OFFSET 17
`define DATA_SINK_FIFO_C2B_CSR_EMPTY 32'h00020000
`define DATA_SINK_FIFO_C2B_CSR_USEDW_OFFSET 0
`define DATA_SINK_FIFO_C2B_CSR_USEDW 32'h000000ff
