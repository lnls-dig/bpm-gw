`define ADDR_WB_FMCPICO1M_4CH_CSR_FMC_STATUS 5'h0
`define WB_FMCPICO1M_4CH_CSR_FMC_STATUS_PRSNT_OFFSET 0
`define WB_FMCPICO1M_4CH_CSR_FMC_STATUS_PRSNT 32'h00000001
`define WB_FMCPICO1M_4CH_CSR_FMC_STATUS_PG_M2C_OFFSET 1
`define WB_FMCPICO1M_4CH_CSR_FMC_STATUS_PG_M2C 32'h00000002
`define ADDR_WB_FMCPICO1M_4CH_CSR_FMC_CTL 5'h4
`define WB_FMCPICO1M_4CH_CSR_FMC_CTL_LED1_OFFSET 0
`define WB_FMCPICO1M_4CH_CSR_FMC_CTL_LED1 32'h00000001
`define WB_FMCPICO1M_4CH_CSR_FMC_CTL_LED2_OFFSET 1
`define WB_FMCPICO1M_4CH_CSR_FMC_CTL_LED2 32'h00000002
`define ADDR_WB_FMCPICO1M_4CH_CSR_RNG_CTL 5'h8
`define WB_FMCPICO1M_4CH_CSR_RNG_CTL_R0_OFFSET 0
`define WB_FMCPICO1M_4CH_CSR_RNG_CTL_R0 32'h00000001
`define WB_FMCPICO1M_4CH_CSR_RNG_CTL_R1_OFFSET 8
`define WB_FMCPICO1M_4CH_CSR_RNG_CTL_R1 32'h00000100
`define WB_FMCPICO1M_4CH_CSR_RNG_CTL_R2_OFFSET 16
`define WB_FMCPICO1M_4CH_CSR_RNG_CTL_R2 32'h00010000
`define WB_FMCPICO1M_4CH_CSR_RNG_CTL_R3_OFFSET 24
`define WB_FMCPICO1M_4CH_CSR_RNG_CTL_R3 32'h01000000
`define ADDR_WB_FMCPICO1M_4CH_CSR_DATA0 5'hc
`define ADDR_WB_FMCPICO1M_4CH_CSR_DATA1 5'h10
`define ADDR_WB_FMCPICO1M_4CH_CSR_DATA2 5'h14
`define ADDR_WB_FMCPICO1M_4CH_CSR_DATA3 5'h18
