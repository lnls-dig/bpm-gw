`define ADDR_FMC150_FLGS_PULSE         5'h0
`define ADDR_FMC150_FLGS_IN            5'h4
`define FMC150_FLGS_IN_SPI_RW_OFFSET 0
`define FMC150_FLGS_IN_SPI_RW 32'h00000001
`define FMC150_FLGS_IN_EXT_CLK_OFFSET 1
`define FMC150_FLGS_IN_EXT_CLK 32'h00000002
`define ADDR_FMC150_ADDR               5'h8
`define ADDR_FMC150_DATA_IN            5'hc
`define ADDR_FMC150_CS                 5'h10
`define FMC150_CS_CDCE72010_OFFSET 0
`define FMC150_CS_CDCE72010 32'h00000001
`define FMC150_CS_ADS62P49_OFFSET 1
`define FMC150_CS_ADS62P49 32'h00000002
`define FMC150_CS_DAC3283_OFFSET 2
`define FMC150_CS_DAC3283 32'h00000004
`define FMC150_CS_AMC7823_OFFSET 3
`define FMC150_CS_AMC7823 32'h00000008
`define ADDR_FMC150_ADC_DLY            5'h14
`define FMC150_ADC_DLY_STR_OFFSET 0
`define FMC150_ADC_DLY_STR 32'h0000001f
`define FMC150_ADC_DLY_CHA_OFFSET 8
`define FMC150_ADC_DLY_CHA 32'h00001f00
`define FMC150_ADC_DLY_CHB_OFFSET 16
`define FMC150_ADC_DLY_CHB 32'h001f0000
`define ADDR_FMC150_DATA_OUT           5'h18
`define ADDR_FMC150_FLGS_OUT           5'h1c
`define FMC150_FLGS_OUT_SPI_BUSY_OFFSET 0
`define FMC150_FLGS_OUT_SPI_BUSY 32'h00000001
`define FMC150_FLGS_OUT_ADC_CLK_LOCKED_OFFSET 1
`define FMC150_FLGS_OUT_ADC_CLK_LOCKED 32'h00000002
