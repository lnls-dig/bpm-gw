`define ADDR_WB_TRIG_IFACE_CH0_CTL     9'h0
`define WB_TRIG_IFACE_CH0_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH0_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH0_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH0_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH0_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH0_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH0_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH0_CTL_TRANSM_COUNT_RST 32'h00000008
`define ADDR_WB_TRIG_IFACE_CH0_CFG     9'h4
`define WB_TRIG_IFACE_CH0_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH0_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH0_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH0_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH0_COUNT   9'h8
`define WB_TRIG_IFACE_CH0_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH0_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH0_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH0_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH1_CTL     9'hc
`define WB_TRIG_IFACE_CH1_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH1_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH1_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH1_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH1_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH1_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH1_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH1_CTL_TRANSM_COUNT_RST 32'h00000008
`define ADDR_WB_TRIG_IFACE_CH1_CFG     9'h10
`define WB_TRIG_IFACE_CH1_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH1_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH1_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH1_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH1_COUNT   9'h14
`define WB_TRIG_IFACE_CH1_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH1_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH1_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH1_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH2_CTL     9'h18
`define WB_TRIG_IFACE_CH2_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH2_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH2_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH2_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH2_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH2_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH2_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH2_CTL_TRANSM_COUNT_RST 32'h00000008
`define ADDR_WB_TRIG_IFACE_CH2_CFG     9'h1c
`define WB_TRIG_IFACE_CH2_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH2_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH2_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH2_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH2_COUNT   9'h20
`define WB_TRIG_IFACE_CH2_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH2_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH2_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH2_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH3_CTL     9'h24
`define WB_TRIG_IFACE_CH3_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH3_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH3_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH3_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH3_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH3_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH3_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH3_CTL_TRANSM_COUNT_RST 32'h00000008
`define ADDR_WB_TRIG_IFACE_CH3_CFG     9'h28
`define WB_TRIG_IFACE_CH3_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH3_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH3_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH3_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH3_COUNT   9'h2c
`define WB_TRIG_IFACE_CH3_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH3_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH3_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH3_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH4_CTL     9'h30
`define WB_TRIG_IFACE_CH4_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH4_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH4_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH4_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH4_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH4_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH4_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH4_CTL_TRANSM_COUNT_RST 32'h00000008
`define ADDR_WB_TRIG_IFACE_CH4_CFG     9'h34
`define WB_TRIG_IFACE_CH4_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH4_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH4_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH4_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH4_COUNT   9'h38
`define WB_TRIG_IFACE_CH4_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH4_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH4_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH4_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH5_CTL     9'h3c
`define WB_TRIG_IFACE_CH5_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH5_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH5_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH5_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH5_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH5_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH5_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH5_CTL_TRANSM_COUNT_RST 32'h00000008
`define ADDR_WB_TRIG_IFACE_CH5_CFG     9'h40
`define WB_TRIG_IFACE_CH5_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH5_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH5_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH5_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH5_COUNT   9'h44
`define WB_TRIG_IFACE_CH5_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH5_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH5_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH5_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH6_CTL     9'h48
`define WB_TRIG_IFACE_CH6_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH6_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH6_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH6_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH6_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH6_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH6_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH6_CTL_TRANSM_COUNT_RST 32'h00000008
`define ADDR_WB_TRIG_IFACE_CH6_CFG     9'h4c
`define WB_TRIG_IFACE_CH6_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH6_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH6_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH6_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH6_COUNT   9'h50
`define WB_TRIG_IFACE_CH6_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH6_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH6_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH6_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH7_CTL     9'h54
`define WB_TRIG_IFACE_CH7_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH7_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH7_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH7_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH7_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH7_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH7_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH7_CTL_TRANSM_COUNT_RST 32'h00000008
`define ADDR_WB_TRIG_IFACE_CH7_CFG     9'h58
`define WB_TRIG_IFACE_CH7_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH7_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH7_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH7_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH7_COUNT   9'h5c
`define WB_TRIG_IFACE_CH7_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH7_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH7_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH7_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH8_CTL     9'h60
`define WB_TRIG_IFACE_CH8_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH8_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH8_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH8_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH8_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH8_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH8_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH8_CTL_TRANSM_COUNT_RST 32'h00000008
`define ADDR_WB_TRIG_IFACE_CH8_CFG     9'h64
`define WB_TRIG_IFACE_CH8_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH8_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH8_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH8_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH8_COUNT   9'h68
`define WB_TRIG_IFACE_CH8_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH8_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH8_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH8_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH9_CTL     9'h6c
`define WB_TRIG_IFACE_CH9_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH9_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH9_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH9_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH9_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH9_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH9_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH9_CTL_TRANSM_COUNT_RST 32'h00000008
`define ADDR_WB_TRIG_IFACE_CH9_CFG     9'h70
`define WB_TRIG_IFACE_CH9_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH9_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH9_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH9_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH9_COUNT   9'h74
`define WB_TRIG_IFACE_CH9_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH9_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH9_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH9_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH10_CTL    9'h78
`define WB_TRIG_IFACE_CH10_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH10_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH10_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH10_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH10_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH10_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH10_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH10_CTL_TRANSM_COUNT_RST 32'h00000008
`define ADDR_WB_TRIG_IFACE_CH10_CFG    9'h7c
`define WB_TRIG_IFACE_CH10_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH10_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH10_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH10_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH10_COUNT  9'h80
`define WB_TRIG_IFACE_CH10_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH10_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH10_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH10_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH11_CTL    9'h84
`define WB_TRIG_IFACE_CH11_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH11_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH11_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH11_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH11_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH11_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH11_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH11_CTL_TRANSM_COUNT_RST 32'h00000008
`define ADDR_WB_TRIG_IFACE_CH11_CFG    9'h88
`define WB_TRIG_IFACE_CH11_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH11_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH11_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH11_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH11_COUNT  9'h8c
`define WB_TRIG_IFACE_CH11_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH11_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH11_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH11_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH12_CTL    9'h90
`define WB_TRIG_IFACE_CH12_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH12_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH12_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH12_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH12_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH12_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH12_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH12_CTL_TRANSM_COUNT_RST 32'h00000008
`define ADDR_WB_TRIG_IFACE_CH12_CFG    9'h94
`define WB_TRIG_IFACE_CH12_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH12_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH12_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH12_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH12_COUNT  9'h98
`define WB_TRIG_IFACE_CH12_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH12_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH12_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH12_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH13_CTL    9'h9c
`define WB_TRIG_IFACE_CH13_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH13_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH13_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH13_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH13_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH13_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH13_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH13_CTL_TRANSM_COUNT_RST 32'h00000008
`define ADDR_WB_TRIG_IFACE_CH13_CFG    9'ha0
`define WB_TRIG_IFACE_CH13_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH13_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH13_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH13_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH13_COUNT  9'ha4
`define WB_TRIG_IFACE_CH13_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH13_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH13_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH13_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH14_CTL    9'ha8
`define WB_TRIG_IFACE_CH14_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH14_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH14_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH14_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH14_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH14_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH14_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH14_CTL_TRANSM_COUNT_RST 32'h00000008
`define ADDR_WB_TRIG_IFACE_CH14_CFG    9'hac
`define WB_TRIG_IFACE_CH14_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH14_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH14_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH14_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH14_COUNT  9'hb0
`define WB_TRIG_IFACE_CH14_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH14_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH14_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH14_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH15_CTL    9'hb4
`define WB_TRIG_IFACE_CH15_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH15_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH15_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH15_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH15_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH15_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH15_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH15_CTL_TRANSM_COUNT_RST 32'h00000008
`define ADDR_WB_TRIG_IFACE_CH15_CFG    9'hb8
`define WB_TRIG_IFACE_CH15_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH15_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH15_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH15_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH15_COUNT  9'hbc
`define WB_TRIG_IFACE_CH15_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH15_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH15_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH15_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH16_CTL    9'hc0
`define WB_TRIG_IFACE_CH16_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH16_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH16_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH16_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH16_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH16_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH16_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH16_CTL_TRANSM_COUNT_RST 32'h00000008
`define ADDR_WB_TRIG_IFACE_CH16_CFG    9'hc4
`define WB_TRIG_IFACE_CH16_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH16_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH16_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH16_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH16_COUNT  9'hc8
`define WB_TRIG_IFACE_CH16_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH16_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH16_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH16_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH17_CTL    9'hcc
`define WB_TRIG_IFACE_CH17_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH17_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH17_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH17_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH17_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH17_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH17_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH17_CTL_TRANSM_COUNT_RST 32'h00000008
`define ADDR_WB_TRIG_IFACE_CH17_CFG    9'hd0
`define WB_TRIG_IFACE_CH17_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH17_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH17_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH17_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH17_COUNT  9'hd4
`define WB_TRIG_IFACE_CH17_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH17_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH17_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH17_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH18_CTL    9'hd8
`define WB_TRIG_IFACE_CH18_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH18_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH18_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH18_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH18_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH18_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH18_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH18_CTL_TRANSM_COUNT_RST 32'h00000008
`define ADDR_WB_TRIG_IFACE_CH18_CFG    9'hdc
`define WB_TRIG_IFACE_CH18_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH18_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH18_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH18_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH18_COUNT  9'he0
`define WB_TRIG_IFACE_CH18_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH18_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH18_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH18_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH19_CTL    9'he4
`define WB_TRIG_IFACE_CH19_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH19_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH19_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH19_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH19_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH19_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH19_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH19_CTL_TRANSM_COUNT_RST 32'h00000008
`define ADDR_WB_TRIG_IFACE_CH19_CFG    9'he8
`define WB_TRIG_IFACE_CH19_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH19_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH19_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH19_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH19_COUNT  9'hec
`define WB_TRIG_IFACE_CH19_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH19_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH19_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH19_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH20_CTL    9'hf0
`define WB_TRIG_IFACE_CH20_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH20_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH20_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH20_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH20_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH20_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH20_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH20_CTL_TRANSM_COUNT_RST 32'h00000008
`define ADDR_WB_TRIG_IFACE_CH20_CFG    9'hf4
`define WB_TRIG_IFACE_CH20_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH20_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH20_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH20_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH20_COUNT  9'hf8
`define WB_TRIG_IFACE_CH20_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH20_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH20_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH20_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH21_CTL    9'hfc
`define WB_TRIG_IFACE_CH21_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH21_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH21_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH21_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH21_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH21_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH21_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH21_CTL_TRANSM_COUNT_RST 32'h00000008
`define ADDR_WB_TRIG_IFACE_CH21_CFG    9'h100
`define WB_TRIG_IFACE_CH21_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH21_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH21_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH21_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH21_COUNT  9'h104
`define WB_TRIG_IFACE_CH21_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH21_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH21_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH21_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH22_CTL    9'h108
`define WB_TRIG_IFACE_CH22_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH22_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH22_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH22_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH22_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH22_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH22_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH22_CTL_TRANSM_COUNT_RST 32'h00000008
`define ADDR_WB_TRIG_IFACE_CH22_CFG    9'h10c
`define WB_TRIG_IFACE_CH22_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH22_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH22_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH22_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH22_COUNT  9'h110
`define WB_TRIG_IFACE_CH22_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH22_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH22_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH22_COUNT_TRANSM 32'hffff0000
`define ADDR_WB_TRIG_IFACE_CH23_CTL    9'h114
`define WB_TRIG_IFACE_CH23_CTL_DIR_OFFSET 0
`define WB_TRIG_IFACE_CH23_CTL_DIR 32'h00000001
`define WB_TRIG_IFACE_CH23_CTL_DIR_POL_OFFSET 1
`define WB_TRIG_IFACE_CH23_CTL_DIR_POL 32'h00000002
`define WB_TRIG_IFACE_CH23_CTL_RCV_COUNT_RST_OFFSET 2
`define WB_TRIG_IFACE_CH23_CTL_RCV_COUNT_RST 32'h00000004
`define WB_TRIG_IFACE_CH23_CTL_TRANSM_COUNT_RST_OFFSET 3
`define WB_TRIG_IFACE_CH23_CTL_TRANSM_COUNT_RST 32'h00000008
`define ADDR_WB_TRIG_IFACE_CH23_CFG    9'h118
`define WB_TRIG_IFACE_CH23_CFG_RCV_LEN_OFFSET 0
`define WB_TRIG_IFACE_CH23_CFG_RCV_LEN 32'h000000ff
`define WB_TRIG_IFACE_CH23_CFG_TRANSM_LEN_OFFSET 8
`define WB_TRIG_IFACE_CH23_CFG_TRANSM_LEN 32'h0000ff00
`define ADDR_WB_TRIG_IFACE_CH23_COUNT  9'h11c
`define WB_TRIG_IFACE_CH23_COUNT_RCV_OFFSET 0
`define WB_TRIG_IFACE_CH23_COUNT_RCV 32'h0000ffff
`define WB_TRIG_IFACE_CH23_COUNT_TRANSM_OFFSET 16
`define WB_TRIG_IFACE_CH23_COUNT_TRANSM 32'hffff0000
